// Generated from: 20250609-202437_binTestAcc9721_seed820279_epochs100_2x1600_b256_lr75_interconnect.pth

module net (
    input  wire [255:0] in,
    output wire [1599:0] out,
    output wire [1269:0] categories
);
    wire [1600:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = in[94]; 
    assign layer_0[1] = ~in[46]; 
    assign layer_0[2] = ~(in[227] | in[243]); 
    assign layer_0[3] = in[234] & ~in[171]; 
    assign layer_0[4] = ~(in[236] ^ in[206]); 
    assign layer_0[5] = ~(in[71] ^ in[41]); 
    assign layer_0[6] = ~in[197]; 
    assign layer_0[7] = in[102] ^ in[115]; 
    assign layer_0[8] = in[148] ^ in[118]; 
    assign layer_0[9] = ~(in[36] | in[21]); 
    assign layer_0[10] = ~in[135] | (in[96] & in[135]); 
    assign layer_0[11] = ~(in[163] ^ in[181]); 
    assign layer_0[12] = in[182] & ~in[53]; 
    assign layer_0[13] = in[55] ^ in[86]; 
    assign layer_0[14] = in[156] | in[163]; 
    assign layer_0[15] = ~in[132]; 
    assign layer_0[16] = in[22] | in[188]; 
    assign layer_0[17] = in[117] | in[55]; 
    assign layer_0[18] = in[157] | in[188]; 
    assign layer_0[19] = ~(in[68] ^ in[191]); 
    assign layer_0[20] = ~in[70] | (in[70] & in[118]); 
    assign layer_0[21] = in[115]; 
    assign layer_0[22] = in[83] | in[167]; 
    assign layer_0[23] = ~(in[218] ^ in[185]); 
    assign layer_0[24] = in[47]; 
    assign layer_0[25] = in[46] | in[51]; 
    assign layer_0[26] = ~(in[155] | in[83]); 
    assign layer_0[27] = in[220] ^ in[189]; 
    assign layer_0[28] = ~(in[60] ^ in[93]); 
    assign layer_0[29] = ~in[40] | (in[164] & in[40]); 
    assign layer_0[30] = in[86] & ~in[135]; 
    assign layer_0[31] = in[65] ^ in[34]; 
    assign layer_0[32] = in[196] & ~in[50]; 
    assign layer_0[33] = in[131] ^ in[117]; 
    assign layer_0[34] = ~in[221] | (in[221] & in[195]); 
    assign layer_0[35] = ~in[135] | (in[219] & in[135]); 
    assign layer_0[36] = ~(in[89] ^ in[75]); 
    assign layer_0[37] = ~in[72] | (in[72] & in[59]); 
    assign layer_0[38] = ~(in[183] ^ in[140]); 
    assign layer_0[39] = ~in[147] | (in[153] & in[147]); 
    assign layer_0[40] = in[132] ^ in[130]; 
    assign layer_0[41] = in[234]; 
    assign layer_0[42] = ~(in[109] | in[107]); 
    assign layer_0[43] = ~(in[165] | in[84]); 
    assign layer_0[44] = in[135] | in[133]; 
    assign layer_0[45] = in[245] & ~in[181]; 
    assign layer_0[46] = in[98] | in[68]; 
    assign layer_0[47] = in[88]; 
    assign layer_0[48] = ~in[170] | (in[170] & in[196]); 
    assign layer_0[49] = ~in[143] | (in[143] & in[109]); 
    assign layer_0[50] = in[242] | in[159]; 
    assign layer_0[51] = ~in[74] | (in[120] & in[74]); 
    assign layer_0[52] = in[139] ^ in[107]; 
    assign layer_0[53] = in[53] ^ in[107]; 
    assign layer_0[54] = ~(in[167] ^ in[83]); 
    assign layer_0[55] = ~in[196]; 
    assign layer_0[56] = in[105] & ~in[78]; 
    assign layer_0[57] = in[120] | in[87]; 
    assign layer_0[58] = in[237] ^ in[205]; 
    assign layer_0[59] = in[172] ^ in[141]; 
    assign layer_0[60] = ~(in[111] | in[79]); 
    assign layer_0[61] = in[177] & ~in[244]; 
    assign layer_0[62] = in[73] & ~in[24]; 
    assign layer_0[63] = in[107] | in[124]; 
    assign layer_0[64] = in[199] ^ in[179]; 
    assign layer_0[65] = in[230] & ~in[10]; 
    assign layer_0[66] = ~in[89] | (in[89] & in[8]); 
    assign layer_0[67] = in[165] ^ in[183]; 
    assign layer_0[68] = ~(in[23] ^ in[214]); 
    assign layer_0[69] = ~in[39] | (in[39] & in[105]); 
    assign layer_0[70] = ~(in[98] ^ in[78]); 
    assign layer_0[71] = ~(in[58] ^ in[89]); 
    assign layer_0[72] = ~(in[22] ^ in[74]); 
    assign layer_0[73] = ~(in[169] | in[154]); 
    assign layer_0[74] = in[56] ^ in[78]; 
    assign layer_0[75] = ~(in[251] ^ in[237]); 
    assign layer_0[76] = ~(in[118] ^ in[173]); 
    assign layer_0[77] = in[164] | in[196]; 
    assign layer_0[78] = ~(in[181] | in[183]); 
    assign layer_0[79] = ~(in[99] ^ in[40]); 
    assign layer_0[80] = ~in[95]; 
    assign layer_0[81] = in[73] ^ in[75]; 
    assign layer_0[82] = in[117] ^ in[130]; 
    assign layer_0[83] = ~(in[120] | in[121]); 
    assign layer_0[84] = ~(in[101] ^ in[67]); 
    assign layer_0[85] = ~in[214] | (in[103] & in[214]); 
    assign layer_0[86] = ~(in[9] ^ in[40]); 
    assign layer_0[87] = ~in[216] | (in[54] & in[216]); 
    assign layer_0[88] = ~(in[199] ^ in[133]); 
    assign layer_0[89] = in[182] & ~in[73]; 
    assign layer_0[90] = ~in[76] | (in[149] & in[76]); 
    assign layer_0[91] = ~in[38]; 
    assign layer_0[92] = in[242] | in[65]; 
    assign layer_0[93] = in[72] & in[102]; 
    assign layer_0[94] = ~(in[195] | in[52]); 
    assign layer_0[95] = in[154] ^ in[20]; 
    assign layer_0[96] = ~(in[179] & in[94]); 
    assign layer_0[97] = ~(in[94] ^ in[166]); 
    assign layer_0[98] = ~(in[19] | in[92]); 
    assign layer_0[99] = ~(in[66] ^ in[38]); 
    assign layer_0[100] = ~(in[110] ^ in[111]); 
    assign layer_0[101] = ~in[23] | (in[23] & in[148]); 
    assign layer_0[102] = in[149] & ~in[106]; 
    assign layer_0[103] = ~(in[183] | in[119]); 
    assign layer_0[104] = ~in[73] | (in[39] & in[73]); 
    assign layer_0[105] = ~(in[99] | in[117]); 
    assign layer_0[106] = ~(in[102] | in[116]); 
    assign layer_0[107] = in[167] | in[150]; 
    assign layer_0[108] = in[165] ^ in[232]; 
    assign layer_0[109] = in[142] ^ in[88]; 
    assign layer_0[110] = in[76] ^ in[72]; 
    assign layer_0[111] = ~in[167] | (in[167] & in[243]); 
    assign layer_0[112] = ~in[170] | (in[170] & in[173]); 
    assign layer_0[113] = ~in[201] | (in[248] & in[201]); 
    assign layer_0[114] = in[137] & ~in[84]; 
    assign layer_0[115] = ~(in[23] ^ in[55]); 
    assign layer_0[116] = in[249] | in[199]; 
    assign layer_0[117] = in[133] & ~in[183]; 
    assign layer_0[118] = ~in[138]; 
    assign layer_0[119] = in[232] | in[216]; 
    assign layer_0[120] = ~in[149] | (in[149] & in[245]); 
    assign layer_0[121] = in[157]; 
    assign layer_0[122] = ~(in[184] ^ in[212]); 
    assign layer_0[123] = in[132] & ~in[81]; 
    assign layer_0[124] = in[130] & in[99]; 
    assign layer_0[125] = ~(in[89] ^ in[42]); 
    assign layer_0[126] = ~in[122] | (in[26] & in[122]); 
    assign layer_0[127] = ~(in[116] ^ in[102]); 
    assign layer_0[128] = in[69] | in[54]; 
    assign layer_0[129] = ~in[211] | (in[105] & in[211]); 
    assign layer_0[130] = in[133] | in[228]; 
    assign layer_0[131] = ~(in[166] | in[183]); 
    assign layer_0[132] = ~(in[71] ^ in[42]); 
    assign layer_0[133] = ~(in[152] ^ in[105]); 
    assign layer_0[134] = ~in[90] | (in[90] & in[116]); 
    assign layer_0[135] = ~(in[30] | in[67]); 
    assign layer_0[136] = ~in[154] | (in[154] & in[200]); 
    assign layer_0[137] = in[205] ^ in[181]; 
    assign layer_0[138] = in[72] ^ in[70]; 
    assign layer_0[139] = in[133] | in[132]; 
    assign layer_0[140] = ~(in[78] ^ in[124]); 
    assign layer_0[141] = ~(in[87] ^ in[101]); 
    assign layer_0[142] = ~(in[214] ^ in[245]); 
    assign layer_0[143] = ~in[72] | (in[47] & in[72]); 
    assign layer_0[144] = in[168] & ~in[37]; 
    assign layer_0[145] = in[70] & ~in[135]; 
    assign layer_0[146] = in[46] | in[29]; 
    assign layer_0[147] = in[106] | in[108]; 
    assign layer_0[148] = in[216] & ~in[131]; 
    assign layer_0[149] = ~(in[90] | in[92]); 
    assign layer_0[150] = ~in[104] | (in[150] & in[104]); 
    assign layer_0[151] = ~(in[214] ^ in[199]); 
    assign layer_0[152] = in[199] ^ in[44]; 
    assign layer_0[153] = ~(in[142] | in[109]); 
    assign layer_0[154] = ~(in[85] ^ in[99]); 
    assign layer_0[155] = ~(in[26] ^ in[45]); 
    assign layer_0[156] = ~in[248] | (in[69] & in[248]); 
    assign layer_0[157] = ~in[129]; 
    assign layer_0[158] = in[82] | in[139]; 
    assign layer_0[159] = in[56] & ~in[214]; 
    assign layer_0[160] = in[59] & in[121]; 
    assign layer_0[161] = in[24] ^ in[79]; 
    assign layer_0[162] = ~in[109]; 
    assign layer_0[163] = ~(in[90] & in[122]); 
    assign layer_0[164] = ~(in[250] | in[90]); 
    assign layer_0[165] = ~(in[191] | in[103]); 
    assign layer_0[166] = ~(in[106] | in[187]); 
    assign layer_0[167] = in[117] ^ in[131]; 
    assign layer_0[168] = ~(in[166] | in[105]); 
    assign layer_0[169] = in[180] & ~in[213]; 
    assign layer_0[170] = ~(in[168] | in[27]); 
    assign layer_0[171] = in[196] | in[228]; 
    assign layer_0[172] = ~(in[156] | in[88]); 
    assign layer_0[173] = in[139] ^ in[140]; 
    assign layer_0[174] = in[179] ^ in[197]; 
    assign layer_0[175] = in[162] | in[121]; 
    assign layer_0[176] = ~(in[72] | in[86]); 
    assign layer_0[177] = in[148] & ~in[151]; 
    assign layer_0[178] = in[229] & ~in[162]; 
    assign layer_0[179] = ~(in[90] & in[74]); 
    assign layer_0[180] = ~in[87] | (in[189] & in[87]); 
    assign layer_0[181] = ~(in[116] ^ in[114]); 
    assign layer_0[182] = ~(in[228] ^ in[182]); 
    assign layer_0[183] = in[167] & ~in[58]; 
    assign layer_0[184] = ~(in[155] | in[53]); 
    assign layer_0[185] = ~(in[127] | in[184]); 
    assign layer_0[186] = in[138] & ~in[195]; 
    assign layer_0[187] = in[73] & in[131]; 
    assign layer_0[188] = ~(in[203] | in[173]); 
    assign layer_0[189] = in[165] ^ in[135]; 
    assign layer_0[190] = ~(in[93] ^ in[107]); 
    assign layer_0[191] = in[103] | in[125]; 
    assign layer_0[192] = in[149] & ~in[167]; 
    assign layer_0[193] = in[156] ^ in[138]; 
    assign layer_0[194] = ~in[229]; 
    assign layer_0[195] = ~(in[251] | in[218]); 
    assign layer_0[196] = ~(in[198] ^ in[244]); 
    assign layer_0[197] = in[136] & in[167]; 
    assign layer_0[198] = ~(in[92] ^ in[73]); 
    assign layer_0[199] = ~(in[26] | in[43]); 
    assign layer_0[200] = ~in[77]; 
    assign layer_0[201] = in[209]; 
    assign layer_0[202] = in[247] & ~in[129]; 
    assign layer_0[203] = in[85] & ~in[211]; 
    assign layer_0[204] = ~(in[41] | in[26]); 
    assign layer_0[205] = ~(in[202] ^ in[233]); 
    assign layer_0[206] = in[51] ^ in[139]; 
    assign layer_0[207] = in[87]; 
    assign layer_0[208] = in[153] & in[122]; 
    assign layer_0[209] = in[38] ^ in[54]; 
    assign layer_0[210] = ~(in[59] ^ in[44]); 
    assign layer_0[211] = ~(in[81] | in[50]); 
    assign layer_0[212] = ~(in[132] ^ in[134]); 
    assign layer_0[213] = in[228] | in[99]; 
    assign layer_0[214] = in[134] & ~in[158]; 
    assign layer_0[215] = ~(in[44] | in[42]); 
    assign layer_0[216] = in[115] | in[102]; 
    assign layer_0[217] = ~(in[124] ^ in[119]); 
    assign layer_0[218] = ~(in[147] | in[11]); 
    assign layer_0[219] = ~(in[212] | in[150]); 
    assign layer_0[220] = ~(in[148] | in[146]); 
    assign layer_0[221] = ~(in[94] | in[88]); 
    assign layer_0[222] = in[88] & ~in[60]; 
    assign layer_0[223] = in[190] | in[171]; 
    assign layer_0[224] = ~(in[92] ^ in[124]); 
    assign layer_0[225] = in[85]; 
    assign layer_0[226] = ~(in[60] | in[180]); 
    assign layer_0[227] = ~in[105] | (in[105] & in[72]); 
    assign layer_0[228] = ~(in[150] | in[168]); 
    assign layer_0[229] = ~(in[154] ^ in[173]); 
    assign layer_0[230] = in[140] | in[123]; 
    assign layer_0[231] = ~(in[137] ^ in[180]); 
    assign layer_0[232] = ~(in[140] | in[155]); 
    assign layer_0[233] = in[69] ^ in[103]; 
    assign layer_0[234] = in[188] | in[54]; 
    assign layer_0[235] = ~in[70] | (in[150] & in[70]); 
    assign layer_0[236] = in[221] | in[204]; 
    assign layer_0[237] = in[55] & ~in[171]; 
    assign layer_0[238] = in[185] & in[54]; 
    assign layer_0[239] = in[90] & ~in[155]; 
    assign layer_0[240] = in[147] ^ in[82]; 
    assign layer_0[241] = in[185] & ~in[221]; 
    assign layer_0[242] = ~in[150] | (in[146] & in[150]); 
    assign layer_0[243] = in[41]; 
    assign layer_0[244] = in[197] | in[198]; 
    assign layer_0[245] = ~(in[118] ^ in[154]); 
    assign layer_0[246] = ~in[179] | (in[179] & in[220]); 
    assign layer_0[247] = in[92] | in[91]; 
    assign layer_0[248] = in[104] & ~in[138]; 
    assign layer_0[249] = in[94] ^ in[151]; 
    assign layer_0[250] = ~(in[172] ^ in[119]); 
    assign layer_0[251] = in[109] ^ in[91]; 
    assign layer_0[252] = in[215]; 
    assign layer_0[253] = ~(in[103] ^ in[153]); 
    assign layer_0[254] = in[148] | in[151]; 
    assign layer_0[255] = in[42] ^ in[52]; 
    assign layer_0[256] = ~in[84] | (in[84] & in[211]); 
    assign layer_0[257] = in[72] ^ in[37]; 
    assign layer_0[258] = in[215] ^ in[212]; 
    assign layer_0[259] = in[21] | in[177]; 
    assign layer_0[260] = in[181] ^ in[229]; 
    assign layer_0[261] = ~in[99] | (in[215] & in[99]); 
    assign layer_0[262] = ~in[148] | (in[148] & in[88]); 
    assign layer_0[263] = ~(in[140] ^ in[122]); 
    assign layer_0[264] = ~in[59] | (in[59] & in[119]); 
    assign layer_0[265] = in[24] & ~in[165]; 
    assign layer_0[266] = in[125] ^ in[108]; 
    assign layer_0[267] = in[98] & ~in[217]; 
    assign layer_0[268] = ~(in[61] ^ in[27]); 
    assign layer_0[269] = ~(in[36] | in[7]); 
    assign layer_0[270] = ~(in[147] | in[130]); 
    assign layer_0[271] = ~(in[180] | in[155]); 
    assign layer_0[272] = ~in[26]; 
    assign layer_0[273] = ~(in[50] | in[81]); 
    assign layer_0[274] = ~(in[138] | in[104]); 
    assign layer_0[275] = in[26] & ~in[59]; 
    assign layer_0[276] = ~(in[166] ^ in[122]); 
    assign layer_0[277] = ~(in[251] ^ in[220]); 
    assign layer_0[278] = ~(in[59] | in[61]); 
    assign layer_0[279] = ~in[129] | (in[129] & in[202]); 
    assign layer_0[280] = in[87] | in[113]; 
    assign layer_0[281] = ~(in[86] ^ in[199]); 
    assign layer_0[282] = ~(in[200] ^ in[115]); 
    assign layer_0[283] = ~in[148] | (in[148] & in[245]); 
    assign layer_0[284] = ~in[137] | (in[137] & in[140]); 
    assign layer_0[285] = in[149] ^ in[119]; 
    assign layer_0[286] = ~in[72] | (in[72] & in[27]); 
    assign layer_0[287] = in[230] ^ in[215]; 
    assign layer_0[288] = in[54] & ~in[8]; 
    assign layer_0[289] = in[162]; 
    assign layer_0[290] = ~(in[36] ^ in[67]); 
    assign layer_0[291] = ~(in[84] | in[98]); 
    assign layer_0[292] = in[30] & ~in[13]; 
    assign layer_0[293] = in[141] ^ in[35]; 
    assign layer_0[294] = in[19] | in[42]; 
    assign layer_0[295] = ~in[105] | (in[105] & in[151]); 
    assign layer_0[296] = in[151] & ~in[81]; 
    assign layer_0[297] = in[165] & ~in[221]; 
    assign layer_0[298] = ~in[183] | (in[231] & in[183]); 
    assign layer_0[299] = ~(in[182] ^ in[78]); 
    assign layer_0[300] = ~(in[233] ^ in[197]); 
    assign layer_0[301] = in[162] ^ in[148]; 
    assign layer_0[302] = ~(in[134] ^ in[103]); 
    assign layer_0[303] = ~in[232] | (in[232] & in[19]); 
    assign layer_0[304] = ~(in[245] | in[244]); 
    assign layer_0[305] = ~in[143] | (in[114] & in[143]); 
    assign layer_0[306] = ~(in[202] | in[82]); 
    assign layer_0[307] = ~(in[103] | in[227]); 
    assign layer_0[308] = in[154]; 
    assign layer_0[309] = ~(in[183] ^ in[180]); 
    assign layer_0[310] = ~in[106] | (in[106] & in[82]); 
    assign layer_0[311] = ~(in[151] ^ in[120]); 
    assign layer_0[312] = in[38]; 
    assign layer_0[313] = ~in[215]; 
    assign layer_0[314] = ~in[40] | (in[21] & in[40]); 
    assign layer_0[315] = in[175] ^ in[195]; 
    assign layer_0[316] = in[131] & ~in[120]; 
    assign layer_0[317] = in[140]; 
    assign layer_0[318] = in[72] ^ in[40]; 
    assign layer_0[319] = ~(in[154] ^ in[122]); 
    assign layer_0[320] = in[163] | in[115]; 
    assign layer_0[321] = ~in[138] | (in[173] & in[138]); 
    assign layer_0[322] = ~(in[58] & in[56]); 
    assign layer_0[323] = in[219] ^ in[172]; 
    assign layer_0[324] = ~(in[247] ^ in[199]); 
    assign layer_0[325] = in[73]; 
    assign layer_0[326] = ~(in[151] & in[182]); 
    assign layer_0[327] = ~in[185] | (in[212] & in[185]); 
    assign layer_0[328] = in[124] | in[142]; 
    assign layer_0[329] = ~(in[153] ^ in[157]); 
    assign layer_0[330] = in[43] & in[40]; 
    assign layer_0[331] = in[87] ^ in[56]; 
    assign layer_0[332] = in[133] & ~in[245]; 
    assign layer_0[333] = in[29] | in[27]; 
    assign layer_0[334] = ~in[151] | (in[230] & in[151]); 
    assign layer_0[335] = ~(in[75] | in[93]); 
    assign layer_0[336] = in[74] | in[75]; 
    assign layer_0[337] = ~(in[116] | in[19]); 
    assign layer_0[338] = in[54] & ~in[123]; 
    assign layer_0[339] = in[233] | in[55]; 
    assign layer_0[340] = ~(in[216] | in[21]); 
    assign layer_0[341] = in[151] ^ in[227]; 
    assign layer_0[342] = in[71] ^ in[101]; 
    assign layer_0[343] = in[231] ^ in[203]; 
    assign layer_0[344] = in[163] & ~in[211]; 
    assign layer_0[345] = in[210] | in[74]; 
    assign layer_0[346] = ~in[155] | (in[22] & in[155]); 
    assign layer_0[347] = in[252] ^ in[41]; 
    assign layer_0[348] = in[67] | in[69]; 
    assign layer_0[349] = ~(in[247] ^ in[168]); 
    assign layer_0[350] = ~(in[75] | in[52]); 
    assign layer_0[351] = ~in[106] | (in[140] & in[106]); 
    assign layer_0[352] = ~(in[198] ^ in[180]); 
    assign layer_0[353] = ~(in[173] | in[188]); 
    assign layer_0[354] = ~(in[226] ^ in[72]); 
    assign layer_0[355] = in[77] ^ in[94]; 
    assign layer_0[356] = ~(in[198] | in[180]); 
    assign layer_0[357] = in[141] ^ in[247]; 
    assign layer_0[358] = in[161] | in[143]; 
    assign layer_0[359] = in[250] ^ in[23]; 
    assign layer_0[360] = in[147] ^ in[166]; 
    assign layer_0[361] = ~(in[117] ^ in[67]); 
    assign layer_0[362] = in[202] ^ in[165]; 
    assign layer_0[363] = in[132] & ~in[38]; 
    assign layer_0[364] = in[183] ^ in[152]; 
    assign layer_0[365] = ~(in[109] ^ in[54]); 
    assign layer_0[366] = ~(in[27] | in[186]); 
    assign layer_0[367] = ~(in[130] | in[100]); 
    assign layer_0[368] = ~(in[195] & in[95]); 
    assign layer_0[369] = ~(in[110] | in[232]); 
    assign layer_0[370] = in[142]; 
    assign layer_0[371] = ~(in[216] & in[217]); 
    assign layer_0[372] = in[140] | in[102]; 
    assign layer_0[373] = ~(in[138] ^ in[169]); 
    assign layer_0[374] = ~in[152] | (in[213] & in[152]); 
    assign layer_0[375] = ~in[250] | (in[204] & in[250]); 
    assign layer_0[376] = ~(in[230] & in[146]); 
    assign layer_0[377] = ~(in[179] | in[182]); 
    assign layer_0[378] = ~(in[103] ^ in[170]); 
    assign layer_0[379] = in[102] & ~in[60]; 
    assign layer_0[380] = in[62]; 
    assign layer_0[381] = in[131] & ~in[249]; 
    assign layer_0[382] = in[119] & ~in[167]; 
    assign layer_0[383] = ~(in[183] ^ in[116]); 
    assign layer_0[384] = ~(in[5] ^ in[151]); 
    assign layer_0[385] = in[102] ^ in[189]; 
    assign layer_0[386] = ~(in[28] ^ in[62]); 
    assign layer_0[387] = in[136]; 
    assign layer_0[388] = in[197] & ~in[46]; 
    assign layer_0[389] = in[120]; 
    assign layer_0[390] = in[91] & ~in[141]; 
    assign layer_0[391] = in[85] ^ in[52]; 
    assign layer_0[392] = ~(in[38] ^ in[70]); 
    assign layer_0[393] = in[65] ^ in[19]; 
    assign layer_0[394] = in[187]; 
    assign layer_0[395] = ~in[251]; 
    assign layer_0[396] = in[119] ^ in[154]; 
    assign layer_0[397] = ~(in[102] ^ in[97]); 
    assign layer_0[398] = in[216] ^ in[169]; 
    assign layer_0[399] = ~(in[29] | in[197]); 
    assign layer_0[400] = in[42] ^ in[73]; 
    assign layer_0[401] = in[199] & ~in[75]; 
    assign layer_0[402] = ~(in[228] ^ in[218]); 
    assign layer_0[403] = ~(in[27] ^ in[57]); 
    assign layer_0[404] = in[117] ^ in[130]; 
    assign layer_0[405] = ~(in[164] ^ in[149]); 
    assign layer_0[406] = ~(in[45] ^ in[94]); 
    assign layer_0[407] = in[251] ^ in[219]; 
    assign layer_0[408] = in[76] & in[138]; 
    assign layer_0[409] = in[5] | in[145]; 
    assign layer_0[410] = in[196] ^ in[186]; 
    assign layer_0[411] = in[170] ^ in[164]; 
    assign layer_0[412] = in[165]; 
    assign layer_0[413] = ~in[142] | (in[138] & in[142]); 
    assign layer_0[414] = in[181] ^ in[229]; 
    assign layer_0[415] = in[107] & ~in[172]; 
    assign layer_0[416] = in[179] & in[131]; 
    assign layer_0[417] = ~in[136] | (in[187] & in[136]); 
    assign layer_0[418] = in[185] ^ in[35]; 
    assign layer_0[419] = ~(in[242] & in[243]); 
    assign layer_0[420] = ~in[168] | (in[186] & in[168]); 
    assign layer_0[421] = ~(in[89] | in[76]); 
    assign layer_0[422] = in[72] & ~in[76]; 
    assign layer_0[423] = in[41] | in[72]; 
    assign layer_0[424] = ~in[198]; 
    assign layer_0[425] = in[243] ^ in[33]; 
    assign layer_0[426] = ~(in[88] ^ in[25]); 
    assign layer_0[427] = ~(in[118] | in[104]); 
    assign layer_0[428] = ~(in[208] | in[4]); 
    assign layer_0[429] = in[169] ^ in[210]; 
    assign layer_0[430] = ~(in[5] | in[207]); 
    assign layer_0[431] = in[155] ^ in[158]; 
    assign layer_0[432] = ~(in[35] | in[74]); 
    assign layer_0[433] = in[55]; 
    assign layer_0[434] = ~in[195]; 
    assign layer_0[435] = ~(in[73] | in[27]); 
    assign layer_0[436] = ~(in[89] ^ in[104]); 
    assign layer_0[437] = in[109]; 
    assign layer_0[438] = in[232] | in[198]; 
    assign layer_0[439] = in[203] ^ in[249]; 
    assign layer_0[440] = ~in[73] | (in[73] & in[195]); 
    assign layer_0[441] = in[20] | in[41]; 
    assign layer_0[442] = in[230] | in[228]; 
    assign layer_0[443] = ~in[54] | (in[54] & in[148]); 
    assign layer_0[444] = in[106] ^ in[73]; 
    assign layer_0[445] = ~(in[139] ^ in[108]); 
    assign layer_0[446] = ~in[171]; 
    assign layer_0[447] = ~(in[62] | in[45]); 
    assign layer_0[448] = ~(in[161] | in[94]); 
    assign layer_0[449] = in[99]; 
    assign layer_0[450] = in[55] & in[168]; 
    assign layer_0[451] = in[107] | in[108]; 
    assign layer_0[452] = ~in[99]; 
    assign layer_0[453] = ~(in[54] | in[170]); 
    assign layer_0[454] = ~(in[231] | in[232]); 
    assign layer_0[455] = in[184] | in[100]; 
    assign layer_0[456] = ~(in[27] ^ in[169]); 
    assign layer_0[457] = ~(in[7] ^ in[21]); 
    assign layer_0[458] = ~(in[102] ^ in[51]); 
    assign layer_0[459] = in[54] ^ in[99]; 
    assign layer_0[460] = ~(in[154] | in[139]); 
    assign layer_0[461] = in[151] ^ in[244]; 
    assign layer_0[462] = ~in[54] | (in[54] & in[110]); 
    assign layer_0[463] = ~in[102] | (in[179] & in[102]); 
    assign layer_0[464] = in[249] ^ in[136]; 
    assign layer_0[465] = in[43] ^ in[74]; 
    assign layer_0[466] = ~in[57] | (in[57] & in[218]); 
    assign layer_0[467] = in[104] ^ in[139]; 
    assign layer_0[468] = ~in[88] | (in[91] & in[88]); 
    assign layer_0[469] = ~(in[103] ^ in[185]); 
    assign layer_0[470] = in[218] & ~in[200]; 
    assign layer_0[471] = ~in[234] | (in[234] & in[170]); 
    assign layer_0[472] = ~(in[75] | in[77]); 
    assign layer_0[473] = ~in[91] | (in[119] & in[91]); 
    assign layer_0[474] = ~(in[70] ^ in[84]); 
    assign layer_0[475] = in[164] ^ in[166]; 
    assign layer_0[476] = in[7] | in[148]; 
    assign layer_0[477] = in[230]; 
    assign layer_0[478] = in[79] | in[34]; 
    assign layer_0[479] = ~(in[8] | in[236]); 
    assign layer_0[480] = in[39] ^ in[71]; 
    assign layer_0[481] = in[181] ^ in[178]; 
    assign layer_0[482] = in[21] ^ in[24]; 
    assign layer_0[483] = in[98] & ~in[85]; 
    assign layer_0[484] = ~(in[99] ^ in[98]); 
    assign layer_0[485] = in[61] ^ in[55]; 
    assign layer_0[486] = in[24] ^ in[70]; 
    assign layer_0[487] = in[210] | in[9]; 
    assign layer_0[488] = in[99] | in[182]; 
    assign layer_0[489] = ~(in[210] | in[74]); 
    assign layer_0[490] = in[108] & ~in[218]; 
    assign layer_0[491] = in[104] | in[146]; 
    assign layer_0[492] = in[85]; 
    assign layer_0[493] = ~(in[186] & in[188]); 
    assign layer_0[494] = ~(in[181] | in[115]); 
    assign layer_0[495] = in[155]; 
    assign layer_0[496] = ~(in[197] ^ in[194]); 
    assign layer_0[497] = in[188] & in[140]; 
    assign layer_0[498] = in[232]; 
    assign layer_0[499] = ~(in[55] ^ in[215]); 
    assign layer_0[500] = in[127] | in[126]; 
    assign layer_0[501] = in[137] & ~in[181]; 
    assign layer_0[502] = in[116] & ~in[206]; 
    assign layer_0[503] = ~in[137] | (in[137] & in[102]); 
    assign layer_0[504] = in[149] | in[246]; 
    assign layer_0[505] = ~in[86] | (in[225] & in[86]); 
    assign layer_0[506] = ~in[43] | (in[90] & in[43]); 
    assign layer_0[507] = ~(in[35] | in[107]); 
    assign layer_0[508] = in[103] ^ in[161]; 
    assign layer_0[509] = in[108] ^ in[110]; 
    assign layer_0[510] = ~(in[146] ^ in[149]); 
    assign layer_0[511] = in[218] | in[186]; 
    assign layer_0[512] = ~(in[116] ^ in[130]); 
    assign layer_0[513] = in[89] & ~in[170]; 
    assign layer_0[514] = in[46] ^ in[79]; 
    assign layer_0[515] = in[195] | in[182]; 
    assign layer_0[516] = in[147]; 
    assign layer_0[517] = in[248] & ~in[38]; 
    assign layer_0[518] = in[10] ^ in[7]; 
    assign layer_0[519] = in[210] | in[84]; 
    assign layer_0[520] = ~in[136] | (in[116] & in[136]); 
    assign layer_0[521] = ~(in[100] ^ in[102]); 
    assign layer_0[522] = in[101] ^ in[115]; 
    assign layer_0[523] = in[103] ^ in[6]; 
    assign layer_0[524] = in[250] ^ in[237]; 
    assign layer_0[525] = ~(in[37] ^ in[185]); 
    assign layer_0[526] = ~(in[184] ^ in[103]); 
    assign layer_0[527] = in[53] & ~in[132]; 
    assign layer_0[528] = in[130] & in[146]; 
    assign layer_0[529] = ~(in[234] ^ in[58]); 
    assign layer_0[530] = in[243] ^ in[212]; 
    assign layer_0[531] = in[78] ^ in[34]; 
    assign layer_0[532] = ~(in[198] | in[197]); 
    assign layer_0[533] = ~(in[93] ^ in[111]); 
    assign layer_0[534] = ~(in[12] ^ in[9]); 
    assign layer_0[535] = ~in[113]; 
    assign layer_0[536] = in[82] ^ in[101]; 
    assign layer_0[537] = ~(in[61] ^ in[92]); 
    assign layer_0[538] = in[46] | in[63]; 
    assign layer_0[539] = ~in[105] | (in[105] & in[166]); 
    assign layer_0[540] = ~(in[37] | in[78]); 
    assign layer_0[541] = ~in[55] | (in[168] & in[55]); 
    assign layer_0[542] = ~(in[66] | in[52]); 
    assign layer_0[543] = in[8] ^ in[242]; 
    assign layer_0[544] = ~(in[136] ^ in[140]); 
    assign layer_0[545] = in[107] | in[35]; 
    assign layer_0[546] = ~in[120] | (in[140] & in[120]); 
    assign layer_0[547] = ~(in[5] | in[110]); 
    assign layer_0[548] = in[149] ^ in[147]; 
    assign layer_0[549] = in[162] & ~in[125]; 
    assign layer_0[550] = ~(in[119] | in[59]); 
    assign layer_0[551] = in[138] ^ in[106]; 
    assign layer_0[552] = ~(in[116] | in[114]); 
    assign layer_0[553] = ~(in[127] ^ in[106]); 
    assign layer_0[554] = ~(in[59] ^ in[107]); 
    assign layer_0[555] = ~(in[69] ^ in[151]); 
    assign layer_0[556] = ~(in[85] ^ in[242]); 
    assign layer_0[557] = in[71] ^ in[68]; 
    assign layer_0[558] = in[120]; 
    assign layer_0[559] = ~(in[87] ^ in[196]); 
    assign layer_0[560] = ~(in[250] | in[173]); 
    assign layer_0[561] = ~(in[26] | in[70]); 
    assign layer_0[562] = ~(in[39] | in[71]); 
    assign layer_0[563] = in[25] | in[40]; 
    assign layer_0[564] = in[30] | in[95]; 
    assign layer_0[565] = ~in[218] | (in[218] & in[171]); 
    assign layer_0[566] = in[46] | in[78]; 
    assign layer_0[567] = ~in[71] | (in[198] & in[71]); 
    assign layer_0[568] = ~(in[56] ^ in[24]); 
    assign layer_0[569] = in[132] | in[231]; 
    assign layer_0[570] = in[40] | in[56]; 
    assign layer_0[571] = ~(in[86] ^ in[100]); 
    assign layer_0[572] = in[57] & ~in[121]; 
    assign layer_0[573] = in[100] ^ in[114]; 
    assign layer_0[574] = in[121] | in[202]; 
    assign layer_0[575] = in[226] | in[37]; 
    assign layer_0[576] = ~(in[223] | in[253]); 
    assign layer_0[577] = ~in[154] | (in[27] & in[154]); 
    assign layer_0[578] = in[243] | in[33]; 
    assign layer_0[579] = in[217] ^ in[214]; 
    assign layer_0[580] = ~in[46]; 
    assign layer_0[581] = in[158] | in[197]; 
    assign layer_0[582] = ~(in[76] ^ in[26]); 
    assign layer_0[583] = in[21] & ~in[53]; 
    assign layer_0[584] = in[249] ^ in[235]; 
    assign layer_0[585] = in[150] | in[252]; 
    assign layer_0[586] = ~(in[99] | in[98]); 
    assign layer_0[587] = in[152] & ~in[157]; 
    assign layer_0[588] = ~in[183] | (in[231] & in[183]); 
    assign layer_0[589] = ~(in[231] ^ in[249]); 
    assign layer_0[590] = in[140] ^ in[115]; 
    assign layer_0[591] = in[40] | in[238]; 
    assign layer_0[592] = in[99] ^ in[68]; 
    assign layer_0[593] = in[118] ^ in[147]; 
    assign layer_0[594] = ~in[139] | (in[139] & in[190]); 
    assign layer_0[595] = ~(in[193] | in[201]); 
    assign layer_0[596] = in[89]; 
    assign layer_0[597] = ~(in[79] | in[43]); 
    assign layer_0[598] = in[187] ^ in[40]; 
    assign layer_0[599] = ~(in[85] ^ in[39]); 
    assign layer_0[600] = in[8] | in[122]; 
    assign layer_0[601] = in[24] ^ in[27]; 
    assign layer_0[602] = ~(in[218] | in[203]); 
    assign layer_0[603] = ~(in[166] ^ in[201]); 
    assign layer_0[604] = in[183] | in[164]; 
    assign layer_0[605] = in[72] & ~in[211]; 
    assign layer_0[606] = ~(in[195] ^ in[38]); 
    assign layer_0[607] = ~(in[139] & in[120]); 
    assign layer_0[608] = ~(in[79] ^ in[114]); 
    assign layer_0[609] = in[146]; 
    assign layer_0[610] = ~(in[152] ^ in[108]); 
    assign layer_0[611] = in[114] ^ in[74]; 
    assign layer_0[612] = in[37] & ~in[68]; 
    assign layer_0[613] = in[74] & ~in[29]; 
    assign layer_0[614] = in[75] | in[126]; 
    assign layer_0[615] = ~(in[40] ^ in[132]); 
    assign layer_0[616] = in[251] ^ in[202]; 
    assign layer_0[617] = in[212] & ~in[242]; 
    assign layer_0[618] = ~(in[63] & in[75]); 
    assign layer_0[619] = ~(in[140] | in[141]); 
    assign layer_0[620] = ~in[125] | (in[125] & in[34]); 
    assign layer_0[621] = in[198] & ~in[243]; 
    assign layer_0[622] = in[88] ^ in[120]; 
    assign layer_0[623] = ~(in[21] | in[132]); 
    assign layer_0[624] = ~(in[20] | in[173]); 
    assign layer_0[625] = ~in[107]; 
    assign layer_0[626] = ~(in[108] | in[171]); 
    assign layer_0[627] = ~in[179] | (in[179] & in[251]); 
    assign layer_0[628] = in[89] ^ in[93]; 
    assign layer_0[629] = ~in[133] | (in[133] & in[67]); 
    assign layer_0[630] = in[121] | in[153]; 
    assign layer_0[631] = ~(in[27] | in[162]); 
    assign layer_0[632] = ~in[184]; 
    assign layer_0[633] = in[146] | in[12]; 
    assign layer_0[634] = in[185] ^ in[69]; 
    assign layer_0[635] = ~(in[90] ^ in[92]); 
    assign layer_0[636] = in[104] & ~in[139]; 
    assign layer_0[637] = in[172] ^ in[140]; 
    assign layer_0[638] = ~(in[108] ^ in[90]); 
    assign layer_0[639] = in[198] | in[195]; 
    assign layer_0[640] = in[116] & ~in[170]; 
    assign layer_0[641] = ~in[138] | (in[138] & in[119]); 
    assign layer_0[642] = in[104] ^ in[74]; 
    assign layer_0[643] = in[94] | in[81]; 
    assign layer_0[644] = in[72] ^ in[74]; 
    assign layer_0[645] = in[183] & ~in[89]; 
    assign layer_0[646] = in[51] ^ in[21]; 
    assign layer_0[647] = in[215] | in[195]; 
    assign layer_0[648] = in[146] ^ in[133]; 
    assign layer_0[649] = ~in[142] | (in[142] & in[154]); 
    assign layer_0[650] = ~in[137] | (in[137] & in[47]); 
    assign layer_0[651] = ~in[23] | (in[85] & in[23]); 
    assign layer_0[652] = in[6] | in[19]; 
    assign layer_0[653] = ~in[177]; 
    assign layer_0[654] = in[65] | in[184]; 
    assign layer_0[655] = in[235] ^ in[189]; 
    assign layer_0[656] = ~(in[246] ^ in[249]); 
    assign layer_0[657] = ~(in[163] | in[139]); 
    assign layer_0[658] = in[170] & ~in[214]; 
    assign layer_0[659] = in[72]; 
    assign layer_0[660] = in[102] ^ in[100]; 
    assign layer_0[661] = in[68] ^ in[249]; 
    assign layer_0[662] = ~in[230] | (in[230] & in[74]); 
    assign layer_0[663] = ~(in[57] ^ in[25]); 
    assign layer_0[664] = in[146] | in[10]; 
    assign layer_0[665] = ~(in[119] ^ in[29]); 
    assign layer_0[666] = ~in[168] | (in[168] & in[149]); 
    assign layer_0[667] = ~(in[243] | in[8]); 
    assign layer_0[668] = in[119] & ~in[204]; 
    assign layer_0[669] = in[105] | in[72]; 
    assign layer_0[670] = ~in[215] | (in[215] & in[155]); 
    assign layer_0[671] = in[248] ^ in[26]; 
    assign layer_0[672] = in[141] | in[143]; 
    assign layer_0[673] = ~(in[116] | in[98]); 
    assign layer_0[674] = ~(in[170] ^ in[156]); 
    assign layer_0[675] = ~(in[254] ^ in[239]); 
    assign layer_0[676] = in[59] ^ in[235]; 
    assign layer_0[677] = ~(in[107] ^ in[138]); 
    assign layer_0[678] = in[182] & ~in[61]; 
    assign layer_0[679] = ~(in[158] ^ in[132]); 
    assign layer_0[680] = ~(in[106] ^ in[167]); 
    assign layer_0[681] = ~(in[252] | in[185]); 
    assign layer_0[682] = ~(in[83] | in[85]); 
    assign layer_0[683] = ~in[107]; 
    assign layer_0[684] = in[195] ^ in[201]; 
    assign layer_0[685] = in[105]; 
    assign layer_0[686] = ~(in[213] ^ in[165]); 
    assign layer_0[687] = ~(in[40] | in[56]); 
    assign layer_0[688] = ~(in[45] ^ in[92]); 
    assign layer_0[689] = ~(in[58] ^ in[90]); 
    assign layer_0[690] = ~(in[88] | in[228]); 
    assign layer_0[691] = in[78] & ~in[131]; 
    assign layer_0[692] = ~(in[69] ^ in[86]); 
    assign layer_0[693] = ~(in[102] | in[100]); 
    assign layer_0[694] = in[117] | in[163]; 
    assign layer_0[695] = in[42] | in[104]; 
    assign layer_0[696] = in[152] ^ in[123]; 
    assign layer_0[697] = ~(in[178] ^ in[120]); 
    assign layer_0[698] = in[153] ^ in[122]; 
    assign layer_0[699] = in[246] ^ in[249]; 
    assign layer_0[700] = ~in[124]; 
    assign layer_0[701] = ~in[232]; 
    assign layer_0[702] = in[227] ^ in[84]; 
    assign layer_0[703] = ~in[171] | (in[171] & in[120]); 
    assign layer_0[704] = in[133] & ~in[42]; 
    assign layer_0[705] = ~(in[63] | in[47]); 
    assign layer_0[706] = ~in[88] | (in[123] & in[88]); 
    assign layer_0[707] = in[245] & ~in[236]; 
    assign layer_0[708] = in[148] ^ in[36]; 
    assign layer_0[709] = ~(in[152] ^ in[95]); 
    assign layer_0[710] = in[57] ^ in[87]; 
    assign layer_0[711] = ~in[203] | (in[203] & in[99]); 
    assign layer_0[712] = ~(in[86] | in[137]); 
    assign layer_0[713] = in[175] ^ in[191]; 
    assign layer_0[714] = ~in[157]; 
    assign layer_0[715] = ~(in[131] | in[114]); 
    assign layer_0[716] = in[97] ^ in[153]; 
    assign layer_0[717] = ~in[29]; 
    assign layer_0[718] = in[167] ^ in[149]; 
    assign layer_0[719] = ~in[197]; 
    assign layer_0[720] = in[52] | in[243]; 
    assign layer_0[721] = ~(in[53] ^ in[55]); 
    assign layer_0[722] = in[99] | in[86]; 
    assign layer_0[723] = ~(in[198] ^ in[201]); 
    assign layer_0[724] = in[120] ^ in[166]; 
    assign layer_0[725] = in[126] ^ in[140]; 
    assign layer_0[726] = in[106]; 
    assign layer_0[727] = ~(in[182] ^ in[152]); 
    assign layer_0[728] = in[104] ^ in[135]; 
    assign layer_0[729] = in[214] & in[214]; 
    assign layer_0[730] = in[156]; 
    assign layer_0[731] = ~(in[199] ^ in[119]); 
    assign layer_0[732] = in[104] | in[57]; 
    assign layer_0[733] = in[253] & in[114]; 
    assign layer_0[734] = ~in[243]; 
    assign layer_0[735] = in[66]; 
    assign layer_0[736] = 1'b0; 
    assign layer_0[737] = in[215] ^ in[247]; 
    assign layer_0[738] = in[92] ^ in[94]; 
    assign layer_0[739] = in[125]; 
    assign layer_0[740] = in[203] | in[186]; 
    assign layer_0[741] = in[164] ^ in[135]; 
    assign layer_0[742] = ~(in[74] ^ in[76]); 
    assign layer_0[743] = in[235] ^ in[38]; 
    assign layer_0[744] = ~(in[188] ^ in[250]); 
    assign layer_0[745] = in[185] | in[107]; 
    assign layer_0[746] = in[55] & ~in[179]; 
    assign layer_0[747] = in[222] ^ in[174]; 
    assign layer_0[748] = ~(in[10] | in[137]); 
    assign layer_0[749] = ~in[133] | (in[133] & in[11]); 
    assign layer_0[750] = in[72] ^ in[41]; 
    assign layer_0[751] = in[197] ^ in[166]; 
    assign layer_0[752] = ~in[120] | (in[120] & in[172]); 
    assign layer_0[753] = ~in[86]; 
    assign layer_0[754] = in[118] & ~in[37]; 
    assign layer_0[755] = in[91] | in[53]; 
    assign layer_0[756] = ~(in[102] ^ in[171]); 
    assign layer_0[757] = ~(in[135] | in[194]); 
    assign layer_0[758] = in[120] ^ in[234]; 
    assign layer_0[759] = ~in[167] | (in[107] & in[167]); 
    assign layer_0[760] = in[24] & ~in[43]; 
    assign layer_0[761] = in[163] & ~in[70]; 
    assign layer_0[762] = in[73] | in[119]; 
    assign layer_0[763] = in[183]; 
    assign layer_0[764] = ~in[219] | (in[149] & in[219]); 
    assign layer_0[765] = ~(in[171] ^ in[35]); 
    assign layer_0[766] = ~(in[142] ^ in[6]); 
    assign layer_0[767] = in[137] & ~in[229]; 
    assign layer_0[768] = ~(in[132] | in[103]); 
    assign layer_0[769] = in[26] ^ in[200]; 
    assign layer_0[770] = ~(in[146] | in[154]); 
    assign layer_0[771] = in[86] & ~in[72]; 
    assign layer_0[772] = ~(in[132] ^ in[166]); 
    assign layer_0[773] = ~(in[148] ^ in[150]); 
    assign layer_0[774] = in[234] | in[203]; 
    assign layer_0[775] = in[57] | in[43]; 
    assign layer_0[776] = in[243] ^ in[67]; 
    assign layer_0[777] = ~in[121] | (in[121] & in[178]); 
    assign layer_0[778] = in[140] | in[157]; 
    assign layer_0[779] = ~(in[230] | in[211]); 
    assign layer_0[780] = ~(in[75] | in[44]); 
    assign layer_0[781] = in[133] ^ in[115]; 
    assign layer_0[782] = in[183] ^ in[229]; 
    assign layer_0[783] = in[21] ^ in[236]; 
    assign layer_0[784] = in[149] | in[147]; 
    assign layer_0[785] = ~in[183] | (in[183] & in[85]); 
    assign layer_0[786] = in[78] ^ in[76]; 
    assign layer_0[787] = in[199] | in[70]; 
    assign layer_0[788] = in[72] ^ in[59]; 
    assign layer_0[789] = in[83] ^ in[202]; 
    assign layer_0[790] = in[117] | in[156]; 
    assign layer_0[791] = ~(in[149] ^ in[185]); 
    assign layer_0[792] = ~in[135] | (in[97] & in[135]); 
    assign layer_0[793] = ~in[106] | (in[71] & in[106]); 
    assign layer_0[794] = ~(in[110] ^ in[109]); 
    assign layer_0[795] = in[213] & ~in[30]; 
    assign layer_0[796] = in[228] ^ in[24]; 
    assign layer_0[797] = in[217] | in[251]; 
    assign layer_0[798] = ~(in[134] ^ in[141]); 
    assign layer_0[799] = ~in[230] | (in[134] & in[230]); 
    assign layer_0[800] = in[180] | in[104]; 
    assign layer_0[801] = in[126] & ~in[130]; 
    assign layer_0[802] = in[119] & ~in[86]; 
    assign layer_0[803] = ~(in[123] | in[36]); 
    assign layer_0[804] = in[197] | in[195]; 
    assign layer_0[805] = ~(in[204] ^ in[13]); 
    assign layer_0[806] = in[185] ^ in[182]; 
    assign layer_0[807] = in[52] ^ in[90]; 
    assign layer_0[808] = in[136] & ~in[182]; 
    assign layer_0[809] = in[88] ^ in[57]; 
    assign layer_0[810] = ~(in[91] ^ in[249]); 
    assign layer_0[811] = in[117] ^ in[162]; 
    assign layer_0[812] = in[162] ^ in[164]; 
    assign layer_0[813] = in[119] | in[134]; 
    assign layer_0[814] = in[211]; 
    assign layer_0[815] = in[105] | in[135]; 
    assign layer_0[816] = in[186] ^ in[69]; 
    assign layer_0[817] = ~(in[122] | in[89]); 
    assign layer_0[818] = in[107] ^ in[244]; 
    assign layer_0[819] = in[118] & ~in[100]; 
    assign layer_0[820] = ~in[117] | (in[117] & in[34]); 
    assign layer_0[821] = in[149] ^ in[148]; 
    assign layer_0[822] = in[79] | in[248]; 
    assign layer_0[823] = in[194] | in[204]; 
    assign layer_0[824] = in[25] | in[195]; 
    assign layer_0[825] = in[57] ^ in[202]; 
    assign layer_0[826] = ~(in[95] ^ in[93]); 
    assign layer_0[827] = in[182] ^ in[164]; 
    assign layer_0[828] = in[148] & ~in[138]; 
    assign layer_0[829] = in[134] & ~in[141]; 
    assign layer_0[830] = ~in[213]; 
    assign layer_0[831] = ~in[247]; 
    assign layer_0[832] = in[98] ^ in[163]; 
    assign layer_0[833] = in[47] ^ in[136]; 
    assign layer_0[834] = in[91] & ~in[8]; 
    assign layer_0[835] = in[118] ^ in[85]; 
    assign layer_0[836] = in[203] ^ in[168]; 
    assign layer_0[837] = ~in[88] | (in[118] & in[88]); 
    assign layer_0[838] = in[136] | in[221]; 
    assign layer_0[839] = in[152] & ~in[38]; 
    assign layer_0[840] = ~in[58] | (in[58] & in[213]); 
    assign layer_0[841] = in[179] | in[180]; 
    assign layer_0[842] = in[205] | in[173]; 
    assign layer_0[843] = ~(in[77] ^ in[75]); 
    assign layer_0[844] = ~(in[250] | in[75]); 
    assign layer_0[845] = in[74]; 
    assign layer_0[846] = ~(in[243] | in[245]); 
    assign layer_0[847] = ~in[243] | (in[243] & in[186]); 
    assign layer_0[848] = in[85] & ~in[215]; 
    assign layer_0[849] = in[58] ^ in[51]; 
    assign layer_0[850] = ~(in[97] ^ in[99]); 
    assign layer_0[851] = in[156] ^ in[197]; 
    assign layer_0[852] = in[45] | in[59]; 
    assign layer_0[853] = in[78]; 
    assign layer_0[854] = ~in[143] | (in[134] & in[143]); 
    assign layer_0[855] = ~(in[85] ^ in[181]); 
    assign layer_0[856] = in[223] ^ in[252]; 
    assign layer_0[857] = in[196] ^ in[187]; 
    assign layer_0[858] = in[105] & ~in[134]; 
    assign layer_0[859] = in[186] ^ in[37]; 
    assign layer_0[860] = in[80] | in[168]; 
    assign layer_0[861] = in[120] ^ in[136]; 
    assign layer_0[862] = ~(in[38] ^ in[70]); 
    assign layer_0[863] = ~(in[179] ^ in[181]); 
    assign layer_0[864] = ~(in[73] & in[28]); 
    assign layer_0[865] = in[167] ^ in[170]; 
    assign layer_0[866] = ~(in[25] ^ in[71]); 
    assign layer_0[867] = ~(in[94] ^ in[46]); 
    assign layer_0[868] = ~(in[132] ^ in[166]); 
    assign layer_0[869] = in[188] | in[183]; 
    assign layer_0[870] = ~(in[164] ^ in[166]); 
    assign layer_0[871] = ~(in[70] ^ in[102]); 
    assign layer_0[872] = in[92] | in[90]; 
    assign layer_0[873] = in[103] & ~in[162]; 
    assign layer_0[874] = ~(in[143] | in[213]); 
    assign layer_0[875] = ~(in[20] | in[78]); 
    assign layer_0[876] = in[196] | in[162]; 
    assign layer_0[877] = ~(in[114] ^ in[100]); 
    assign layer_0[878] = in[145]; 
    assign layer_0[879] = in[154] & ~in[197]; 
    assign layer_0[880] = in[149] ^ in[179]; 
    assign layer_0[881] = ~(in[26] ^ in[57]); 
    assign layer_0[882] = ~(in[19] | in[211]); 
    assign layer_0[883] = in[83] | in[98]; 
    assign layer_0[884] = in[184] ^ in[149]; 
    assign layer_0[885] = in[134] ^ in[165]; 
    assign layer_0[886] = in[170] ^ in[139]; 
    assign layer_0[887] = ~in[119] | (in[119] & in[201]); 
    assign layer_0[888] = ~(in[69] | in[107]); 
    assign layer_0[889] = ~(in[163] ^ in[165]); 
    assign layer_0[890] = in[137] ^ in[117]; 
    assign layer_0[891] = ~(in[12] | in[11]); 
    assign layer_0[892] = ~(in[25] | in[95]); 
    assign layer_0[893] = in[82] & ~in[230]; 
    assign layer_0[894] = in[132] ^ in[158]; 
    assign layer_0[895] = in[89] ^ in[107]; 
    assign layer_0[896] = ~(in[151] | in[136]); 
    assign layer_0[897] = ~(in[130] | in[171]); 
    assign layer_0[898] = ~(in[137] | in[9]); 
    assign layer_0[899] = in[94]; 
    assign layer_0[900] = ~(in[139] ^ in[181]); 
    assign layer_0[901] = in[182] & ~in[172]; 
    assign layer_0[902] = ~(in[220] | in[203]); 
    assign layer_0[903] = ~(in[143] | in[196]); 
    assign layer_0[904] = in[229] ^ in[214]; 
    assign layer_0[905] = in[22] ^ in[41]; 
    assign layer_0[906] = in[204] ^ in[173]; 
    assign layer_0[907] = in[129] & ~in[44]; 
    assign layer_0[908] = in[82] ^ in[52]; 
    assign layer_0[909] = in[57] & ~in[139]; 
    assign layer_0[910] = ~(in[214] ^ in[245]); 
    assign layer_0[911] = ~(in[134] ^ in[126]); 
    assign layer_0[912] = in[103] & in[87]; 
    assign layer_0[913] = in[231] ^ in[92]; 
    assign layer_0[914] = ~(in[9] ^ in[159]); 
    assign layer_0[915] = in[209] | in[205]; 
    assign layer_0[916] = ~(in[179] | in[210]); 
    assign layer_0[917] = in[211] | in[213]; 
    assign layer_0[918] = ~in[131]; 
    assign layer_0[919] = ~in[216] | (in[216] & in[40]); 
    assign layer_0[920] = in[197] ^ in[150]; 
    assign layer_0[921] = ~(in[115] ^ in[113]); 
    assign layer_0[922] = in[149] ^ in[147]; 
    assign layer_0[923] = in[10] | in[211]; 
    assign layer_0[924] = in[138] | in[249]; 
    assign layer_0[925] = ~(in[76] | in[83]); 
    assign layer_0[926] = in[101] ^ in[171]; 
    assign layer_0[927] = ~(in[251] | in[87]); 
    assign layer_0[928] = in[107] ^ in[125]; 
    assign layer_0[929] = in[27] ^ in[60]; 
    assign layer_0[930] = in[124] & in[59]; 
    assign layer_0[931] = in[137] & ~in[187]; 
    assign layer_0[932] = in[164] & ~in[234]; 
    assign layer_0[933] = in[92] ^ in[55]; 
    assign layer_0[934] = in[147] & ~in[119]; 
    assign layer_0[935] = in[136] & ~in[233]; 
    assign layer_0[936] = in[133] ^ in[131]; 
    assign layer_0[937] = ~(in[105] & in[167]); 
    assign layer_0[938] = ~(in[76] | in[104]); 
    assign layer_0[939] = ~in[122]; 
    assign layer_0[940] = in[142] & ~in[153]; 
    assign layer_0[941] = ~(in[195] ^ in[204]); 
    assign layer_0[942] = ~in[88] | (in[88] & in[37]); 
    assign layer_0[943] = in[44] & ~in[141]; 
    assign layer_0[944] = ~(in[112] | in[37]); 
    assign layer_0[945] = in[241] | in[12]; 
    assign layer_0[946] = in[203] ^ in[251]; 
    assign layer_0[947] = in[231] & ~in[104]; 
    assign layer_0[948] = in[39] | in[86]; 
    assign layer_0[949] = ~(in[229] ^ in[196]); 
    assign layer_0[950] = in[103] ^ in[169]; 
    assign layer_0[951] = ~(in[212] ^ in[245]); 
    assign layer_0[952] = in[122] | in[124]; 
    assign layer_0[953] = in[155] | in[54]; 
    assign layer_0[954] = in[29] & ~in[91]; 
    assign layer_0[955] = ~(in[29] ^ in[73]); 
    assign layer_0[956] = in[126]; 
    assign layer_0[957] = in[42] ^ in[52]; 
    assign layer_0[958] = in[112] ^ in[241]; 
    assign layer_0[959] = ~(in[88] ^ in[68]); 
    assign layer_0[960] = in[168] & ~in[123]; 
    assign layer_0[961] = in[134] & ~in[100]; 
    assign layer_0[962] = in[172] | in[155]; 
    assign layer_0[963] = in[45] & ~in[54]; 
    assign layer_0[964] = ~(in[165] | in[148]); 
    assign layer_0[965] = ~(in[228] ^ in[213]); 
    assign layer_0[966] = in[63] ^ in[30]; 
    assign layer_0[967] = ~(in[217] ^ in[28]); 
    assign layer_0[968] = ~in[168] | (in[92] & in[168]); 
    assign layer_0[969] = in[93] ^ in[91]; 
    assign layer_0[970] = ~in[92] | (in[120] & in[92]); 
    assign layer_0[971] = in[86] ^ in[221]; 
    assign layer_0[972] = in[218] & ~in[125]; 
    assign layer_0[973] = in[167] | in[98]; 
    assign layer_0[974] = ~in[153] | (in[195] & in[153]); 
    assign layer_0[975] = ~(in[9] | in[72]); 
    assign layer_0[976] = in[106] ^ in[110]; 
    assign layer_0[977] = ~in[138] | (in[138] & in[157]); 
    assign layer_0[978] = ~(in[193] | in[142]); 
    assign layer_0[979] = ~in[172] | (in[172] & in[170]); 
    assign layer_0[980] = ~in[136]; 
    assign layer_0[981] = ~(in[228] | in[45]); 
    assign layer_0[982] = ~in[214] | (in[214] & in[105]); 
    assign layer_0[983] = in[133] ^ in[147]; 
    assign layer_0[984] = in[119] & ~in[71]; 
    assign layer_0[985] = in[189] ^ in[196]; 
    assign layer_0[986] = in[86]; 
    assign layer_0[987] = in[149]; 
    assign layer_0[988] = in[56] ^ in[103]; 
    assign layer_0[989] = in[93] ^ in[91]; 
    assign layer_0[990] = in[10] & ~in[210]; 
    assign layer_0[991] = in[90] & ~in[141]; 
    assign layer_0[992] = in[75] & ~in[122]; 
    assign layer_0[993] = ~(in[119] ^ in[139]); 
    assign layer_0[994] = ~(in[182] ^ in[180]); 
    assign layer_0[995] = ~(in[67] ^ in[155]); 
    assign layer_0[996] = ~(in[76] ^ in[25]); 
    assign layer_0[997] = ~(in[181] | in[99]); 
    assign layer_0[998] = ~(in[91] | in[183]); 
    assign layer_0[999] = in[181] ^ in[199]; 
    assign layer_0[1000] = ~(in[121] ^ in[171]); 
    assign layer_0[1001] = in[215] & ~in[166]; 
    assign layer_0[1002] = in[113] | in[116]; 
    assign layer_0[1003] = ~(in[99] ^ in[85]); 
    assign layer_0[1004] = in[115] | in[52]; 
    assign layer_0[1005] = in[211] ^ in[189]; 
    assign layer_0[1006] = in[218] & ~in[100]; 
    assign layer_0[1007] = in[86] ^ in[103]; 
    assign layer_0[1008] = ~in[183] | (in[183] & in[186]); 
    assign layer_0[1009] = in[170] ^ in[105]; 
    assign layer_0[1010] = in[88] ^ in[103]; 
    assign layer_0[1011] = ~(in[250] & in[199]); 
    assign layer_0[1012] = in[62] | in[74]; 
    assign layer_0[1013] = ~in[134] | (in[134] & in[218]); 
    assign layer_0[1014] = in[199] & ~in[92]; 
    assign layer_0[1015] = ~(in[213] ^ in[194]); 
    assign layer_0[1016] = in[136] ^ in[104]; 
    assign layer_0[1017] = in[235] ^ in[35]; 
    assign layer_0[1018] = ~(in[69] ^ in[72]); 
    assign layer_0[1019] = in[88] ^ in[101]; 
    assign layer_0[1020] = in[251] & ~in[32]; 
    assign layer_0[1021] = ~in[143]; 
    assign layer_0[1022] = ~(in[107] | in[155]); 
    assign layer_0[1023] = in[251] | in[152]; 
    assign layer_0[1024] = in[105] | in[235]; 
    assign layer_0[1025] = ~(in[219] ^ in[183]); 
    assign layer_0[1026] = ~(in[172] ^ in[138]); 
    assign layer_0[1027] = in[220]; 
    assign layer_0[1028] = ~(in[10] | in[63]); 
    assign layer_0[1029] = ~(in[152] ^ in[199]); 
    assign layer_0[1030] = ~in[134]; 
    assign layer_0[1031] = ~(in[146] | in[139]); 
    assign layer_0[1032] = ~(in[187] | in[186]); 
    assign layer_0[1033] = ~in[170]; 
    assign layer_0[1034] = ~in[184] | (in[61] & in[184]); 
    assign layer_0[1035] = ~(in[163] | in[133]); 
    assign layer_0[1036] = ~in[173]; 
    assign layer_0[1037] = ~(in[58] ^ in[89]); 
    assign layer_0[1038] = ~(in[83] ^ in[52]); 
    assign layer_0[1039] = ~(in[130] | in[163]); 
    assign layer_0[1040] = ~(in[200] | in[182]); 
    assign layer_0[1041] = ~in[213] | (in[213] & in[19]); 
    assign layer_0[1042] = ~(in[62] | in[27]); 
    assign layer_0[1043] = ~(in[135] ^ in[165]); 
    assign layer_0[1044] = in[45]; 
    assign layer_0[1045] = ~in[168] | (in[168] & in[148]); 
    assign layer_0[1046] = in[220] ^ in[181]; 
    assign layer_0[1047] = ~in[87] | (in[52] & in[87]); 
    assign layer_0[1048] = ~(in[120] & in[76]); 
    assign layer_0[1049] = ~(in[38] | in[7]); 
    assign layer_0[1050] = in[146] ^ in[163]; 
    assign layer_0[1051] = ~(in[83] | in[68]); 
    assign layer_0[1052] = in[37] | in[135]; 
    assign layer_0[1053] = in[182] ^ in[151]; 
    assign layer_0[1054] = in[235] | in[106]; 
    assign layer_0[1055] = in[244] & ~in[232]; 
    assign layer_0[1056] = ~(in[30] | in[12]); 
    assign layer_0[1057] = ~in[153] | (in[125] & in[153]); 
    assign layer_0[1058] = ~(in[97] ^ in[99]); 
    assign layer_0[1059] = ~(in[25] ^ in[56]); 
    assign layer_0[1060] = ~(in[149] ^ in[131]); 
    assign layer_0[1061] = in[206] ^ in[85]; 
    assign layer_0[1062] = ~in[88] | (in[77] & in[88]); 
    assign layer_0[1063] = in[111] ^ in[109]; 
    assign layer_0[1064] = in[210] | in[51]; 
    assign layer_0[1065] = in[168] & ~in[126]; 
    assign layer_0[1066] = ~(in[147] ^ in[218]); 
    assign layer_0[1067] = in[87] & ~in[36]; 
    assign layer_0[1068] = ~(in[115] ^ in[129]); 
    assign layer_0[1069] = in[30] ^ in[115]; 
    assign layer_0[1070] = in[71] ^ in[90]; 
    assign layer_0[1071] = ~(in[167] & in[198]); 
    assign layer_0[1072] = in[172] ^ in[165]; 
    assign layer_0[1073] = in[135] ^ in[186]; 
    assign layer_0[1074] = in[150] & in[180]; 
    assign layer_0[1075] = in[140] | in[156]; 
    assign layer_0[1076] = ~(in[189] ^ in[187]); 
    assign layer_0[1077] = ~(in[116] ^ in[102]); 
    assign layer_0[1078] = in[103] ^ in[185]; 
    assign layer_0[1079] = in[181] ^ in[164]; 
    assign layer_0[1080] = ~(in[147] ^ in[171]); 
    assign layer_0[1081] = in[148] ^ in[147]; 
    assign layer_0[1082] = in[168] & in[184]; 
    assign layer_0[1083] = ~(in[165] | in[163]); 
    assign layer_0[1084] = in[100] ^ in[114]; 
    assign layer_0[1085] = in[108] & ~in[249]; 
    assign layer_0[1086] = in[230] ^ in[236]; 
    assign layer_0[1087] = in[165] ^ in[182]; 
    assign layer_0[1088] = ~(in[59] | in[58]); 
    assign layer_0[1089] = in[21] | in[159]; 
    assign layer_0[1090] = in[89] | in[92]; 
    assign layer_0[1091] = ~(in[106] | in[116]); 
    assign layer_0[1092] = ~(in[148] | in[146]); 
    assign layer_0[1093] = ~in[68] | (in[211] & in[68]); 
    assign layer_0[1094] = in[73] & ~in[70]; 
    assign layer_0[1095] = ~(in[118] & in[151]); 
    assign layer_0[1096] = ~in[186] | (in[228] & in[186]); 
    assign layer_0[1097] = in[214] & ~in[227]; 
    assign layer_0[1098] = ~(in[130] ^ in[57]); 
    assign layer_0[1099] = ~(in[217] | in[234]); 
    assign layer_0[1100] = ~(in[52] | in[81]); 
    assign layer_0[1101] = ~(in[140] ^ in[121]); 
    assign layer_0[1102] = in[250] ^ in[84]; 
    assign layer_0[1103] = in[40] | in[132]; 
    assign layer_0[1104] = 1'b1; 
    assign layer_0[1105] = ~(in[149] ^ in[42]); 
    assign layer_0[1106] = ~in[39]; 
    assign layer_0[1107] = ~(in[77] | in[230]); 
    assign layer_0[1108] = ~(in[52] | in[24]); 
    assign layer_0[1109] = in[43] ^ in[76]; 
    assign layer_0[1110] = in[97] | in[98]; 
    assign layer_0[1111] = ~in[57] | (in[184] & in[57]); 
    assign layer_0[1112] = ~(in[141] & in[201]); 
    assign layer_0[1113] = ~in[170] | (in[24] & in[170]); 
    assign layer_0[1114] = in[211] | in[196]; 
    assign layer_0[1115] = ~(in[41] ^ in[43]); 
    assign layer_0[1116] = in[142] | in[29]; 
    assign layer_0[1117] = ~(in[166] ^ in[119]); 
    assign layer_0[1118] = ~in[87] | (in[87] & in[68]); 
    assign layer_0[1119] = ~(in[20] ^ in[7]); 
    assign layer_0[1120] = ~(in[45] | in[76]); 
    assign layer_0[1121] = in[171] & ~in[37]; 
    assign layer_0[1122] = in[216] & ~in[141]; 
    assign layer_0[1123] = ~(in[125] | in[39]); 
    assign layer_0[1124] = ~(in[179] | in[20]); 
    assign layer_0[1125] = ~(in[94] | in[53]); 
    assign layer_0[1126] = ~(in[89] | in[53]); 
    assign layer_0[1127] = ~in[86] | (in[72] & in[86]); 
    assign layer_0[1128] = in[113] ^ in[24]; 
    assign layer_0[1129] = in[5] | in[211]; 
    assign layer_0[1130] = ~in[205] | (in[203] & in[205]); 
    assign layer_0[1131] = in[28] ^ in[142]; 
    assign layer_0[1132] = in[141] & ~in[41]; 
    assign layer_0[1133] = in[216] | in[201]; 
    assign layer_0[1134] = ~(in[164] | in[182]); 
    assign layer_0[1135] = ~in[201] | (in[61] & in[201]); 
    assign layer_0[1136] = ~in[214] | (in[214] & in[75]); 
    assign layer_0[1137] = ~in[45] | (in[45] & in[109]); 
    assign layer_0[1138] = ~(in[26] ^ in[28]); 
    assign layer_0[1139] = ~(in[243] | in[164]); 
    assign layer_0[1140] = ~in[40] | (in[40] & in[237]); 
    assign layer_0[1141] = in[44] ^ in[76]; 
    assign layer_0[1142] = in[89] | in[81]; 
    assign layer_0[1143] = in[229] ^ in[56]; 
    assign layer_0[1144] = in[189] | in[189]; 
    assign layer_0[1145] = ~(in[175] ^ in[88]); 
    assign layer_0[1146] = in[245]; 
    assign layer_0[1147] = in[186] ^ in[234]; 
    assign layer_0[1148] = ~(in[57] ^ in[188]); 
    assign layer_0[1149] = ~in[83] | (in[150] & in[83]); 
    assign layer_0[1150] = ~(in[233] ^ in[180]); 
    assign layer_0[1151] = in[107] | in[235]; 
    assign layer_0[1152] = in[126]; 
    assign layer_0[1153] = in[101] ^ in[170]; 
    assign layer_0[1154] = ~in[124]; 
    assign layer_0[1155] = in[98] ^ in[85]; 
    assign layer_0[1156] = ~(in[91] | in[77]); 
    assign layer_0[1157] = in[126] ^ in[154]; 
    assign layer_0[1158] = ~(in[121] ^ in[99]); 
    assign layer_0[1159] = in[83] ^ in[69]; 
    assign layer_0[1160] = ~(in[71] | in[88]); 
    assign layer_0[1161] = in[60] | in[78]; 
    assign layer_0[1162] = in[147] ^ in[90]; 
    assign layer_0[1163] = ~(in[75] ^ in[73]); 
    assign layer_0[1164] = ~(in[86] | in[99]); 
    assign layer_0[1165] = ~(in[164] ^ in[134]); 
    assign layer_0[1166] = in[247] ^ in[216]; 
    assign layer_0[1167] = in[57] ^ in[59]; 
    assign layer_0[1168] = ~in[117] | (in[117] & in[93]); 
    assign layer_0[1169] = ~in[213]; 
    assign layer_0[1170] = in[203] ^ in[180]; 
    assign layer_0[1171] = in[182] & ~in[232]; 
    assign layer_0[1172] = ~in[152] | (in[146] & in[152]); 
    assign layer_0[1173] = in[197] & ~in[52]; 
    assign layer_0[1174] = in[113] | in[98]; 
    assign layer_0[1175] = ~(in[190] ^ in[221]); 
    assign layer_0[1176] = in[111] ^ in[109]; 
    assign layer_0[1177] = ~(in[229] | in[247]); 
    assign layer_0[1178] = in[204] & ~in[234]; 
    assign layer_0[1179] = in[104] & ~in[78]; 
    assign layer_0[1180] = ~(in[101] ^ in[202]); 
    assign layer_0[1181] = ~(in[244] | in[203]); 
    assign layer_0[1182] = ~in[131]; 
    assign layer_0[1183] = ~(in[76] | in[244]); 
    assign layer_0[1184] = ~(in[59] & in[90]); 
    assign layer_0[1185] = in[162] ^ in[164]; 
    assign layer_0[1186] = in[101] | in[250]; 
    assign layer_0[1187] = in[150] ^ in[84]; 
    assign layer_0[1188] = ~(in[125] ^ in[93]); 
    assign layer_0[1189] = ~in[245] | (in[245] & in[212]); 
    assign layer_0[1190] = ~(in[120] & in[138]); 
    assign layer_0[1191] = in[23] | in[190]; 
    assign layer_0[1192] = ~(in[87] ^ in[242]); 
    assign layer_0[1193] = in[59] ^ in[89]; 
    assign layer_0[1194] = in[114] | in[169]; 
    assign layer_0[1195] = ~(in[91] | in[108]); 
    assign layer_0[1196] = in[177] ^ in[151]; 
    assign layer_0[1197] = in[5] | in[122]; 
    assign layer_0[1198] = in[107] | in[52]; 
    assign layer_0[1199] = ~(in[253] | in[82]); 
    assign layer_0[1200] = ~(in[19] | in[89]); 
    assign layer_0[1201] = ~in[104] | (in[61] & in[104]); 
    assign layer_0[1202] = ~(in[25] & in[172]); 
    assign layer_0[1203] = ~(in[121] ^ in[152]); 
    assign layer_0[1204] = in[161]; 
    assign layer_0[1205] = in[93]; 
    assign layer_0[1206] = in[56] | in[55]; 
    assign layer_0[1207] = ~(in[245] | in[213]); 
    assign layer_0[1208] = ~in[116] | (in[233] & in[116]); 
    assign layer_0[1209] = ~in[151] | (in[163] & in[151]); 
    assign layer_0[1210] = in[211] | in[199]; 
    assign layer_0[1211] = in[180] ^ in[149]; 
    assign layer_0[1212] = in[69] & ~in[23]; 
    assign layer_0[1213] = ~(in[154] | in[94]); 
    assign layer_0[1214] = ~(in[51] | in[221]); 
    assign layer_0[1215] = ~(in[104] | in[11]); 
    assign layer_0[1216] = in[156] | in[38]; 
    assign layer_0[1217] = in[123] ^ in[63]; 
    assign layer_0[1218] = in[237] | in[221]; 
    assign layer_0[1219] = in[177] | in[243]; 
    assign layer_0[1220] = in[167] & ~in[46]; 
    assign layer_0[1221] = in[130] | in[132]; 
    assign layer_0[1222] = ~(in[42] ^ in[68]); 
    assign layer_0[1223] = in[218] & ~in[181]; 
    assign layer_0[1224] = ~(in[58] ^ in[171]); 
    assign layer_0[1225] = ~(in[147] | in[193]); 
    assign layer_0[1226] = ~in[95]; 
    assign layer_0[1227] = ~(in[177] ^ in[168]); 
    assign layer_0[1228] = in[74] & ~in[62]; 
    assign layer_0[1229] = ~(in[104] ^ in[140]); 
    assign layer_0[1230] = ~(in[130] ^ in[117]); 
    assign layer_0[1231] = ~(in[165] | in[230]); 
    assign layer_0[1232] = ~(in[146] ^ in[121]); 
    assign layer_0[1233] = in[100] & ~in[183]; 
    assign layer_0[1234] = ~in[230] | (in[230] & in[121]); 
    assign layer_0[1235] = ~(in[69] ^ in[23]); 
    assign layer_0[1236] = ~(in[172] ^ in[89]); 
    assign layer_0[1237] = in[153] & in[90]; 
    assign layer_0[1238] = in[84] & ~in[86]; 
    assign layer_0[1239] = ~(in[93] & in[90]); 
    assign layer_0[1240] = in[198] ^ in[162]; 
    assign layer_0[1241] = in[167] ^ in[136]; 
    assign layer_0[1242] = in[59] ^ in[27]; 
    assign layer_0[1243] = in[89] ^ in[58]; 
    assign layer_0[1244] = ~(in[194] | in[205]); 
    assign layer_0[1245] = in[249] ^ in[201]; 
    assign layer_0[1246] = in[166]; 
    assign layer_0[1247] = in[247] | in[206]; 
    assign layer_0[1248] = in[210] ^ in[242]; 
    assign layer_0[1249] = in[90] ^ in[108]; 
    assign layer_0[1250] = ~(in[181] | in[183]); 
    assign layer_0[1251] = ~(in[243] ^ in[114]); 
    assign layer_0[1252] = ~in[215] | (in[168] & in[215]); 
    assign layer_0[1253] = in[230]; 
    assign layer_0[1254] = ~(in[235] | in[23]); 
    assign layer_0[1255] = ~in[132] | (in[42] & in[132]); 
    assign layer_0[1256] = ~(in[105] | in[210]); 
    assign layer_0[1257] = in[106] | in[22]; 
    assign layer_0[1258] = ~in[158]; 
    assign layer_0[1259] = ~(in[182] ^ in[155]); 
    assign layer_0[1260] = ~(in[212] | in[5]); 
    assign layer_0[1261] = in[156] ^ in[52]; 
    assign layer_0[1262] = ~(in[133] | in[110]); 
    assign layer_0[1263] = ~in[242]; 
    assign layer_0[1264] = ~(in[104] ^ in[211]); 
    assign layer_0[1265] = ~(in[219] ^ in[201]); 
    assign layer_0[1266] = ~(in[88] ^ in[211]); 
    assign layer_0[1267] = ~(in[206] ^ in[196]); 
    assign layer_0[1268] = in[87] ^ in[90]; 
    assign layer_0[1269] = in[92] | in[146]; 
    assign layer_0[1270] = in[116] & in[131]; 
    assign layer_0[1271] = ~(in[217] | in[233]); 
    assign layer_0[1272] = in[136] & ~in[200]; 
    assign layer_0[1273] = in[168] ^ in[121]; 
    assign layer_0[1274] = ~in[103] | (in[103] & in[35]); 
    assign layer_0[1275] = in[139] & ~in[177]; 
    assign layer_0[1276] = ~(in[206] ^ in[237]); 
    assign layer_0[1277] = ~(in[203] | in[227]); 
    assign layer_0[1278] = ~(in[130] ^ in[116]); 
    assign layer_0[1279] = in[168] & ~in[194]; 
    assign layer_0[1280] = in[103] | in[60]; 
    assign layer_0[1281] = in[138] & ~in[26]; 
    assign layer_0[1282] = ~(in[170] | in[109]); 
    assign layer_0[1283] = ~(in[167] ^ in[165]); 
    assign layer_0[1284] = ~(in[197] ^ in[83]); 
    assign layer_0[1285] = ~in[163] | (in[232] & in[163]); 
    assign layer_0[1286] = ~in[6]; 
    assign layer_0[1287] = in[212] & in[203]; 
    assign layer_0[1288] = ~(in[134] ^ in[9]); 
    assign layer_0[1289] = ~(in[195] ^ in[199]); 
    assign layer_0[1290] = ~(in[56] ^ in[25]); 
    assign layer_0[1291] = ~(in[193] ^ in[174]); 
    assign layer_0[1292] = ~in[170] | (in[170] & in[235]); 
    assign layer_0[1293] = ~in[59] | (in[59] & in[232]); 
    assign layer_0[1294] = ~(in[22] ^ in[36]); 
    assign layer_0[1295] = in[178] ^ in[210]; 
    assign layer_0[1296] = in[178] | in[197]; 
    assign layer_0[1297] = in[71] ^ in[39]; 
    assign layer_0[1298] = ~(in[204] ^ in[154]); 
    assign layer_0[1299] = in[87] | in[101]; 
    assign layer_0[1300] = ~(in[126] ^ in[90]); 
    assign layer_0[1301] = ~(in[85] ^ in[244]); 
    assign layer_0[1302] = in[106] & ~in[219]; 
    assign layer_0[1303] = in[199] & ~in[181]; 
    assign layer_0[1304] = ~(in[198] ^ in[243]); 
    assign layer_0[1305] = ~(in[84] ^ in[98]); 
    assign layer_0[1306] = ~(in[114] | in[132]); 
    assign layer_0[1307] = ~(in[237] | in[153]); 
    assign layer_0[1308] = ~(in[150] & in[170]); 
    assign layer_0[1309] = in[79] & ~in[117]; 
    assign layer_0[1310] = ~(in[139] | in[125]); 
    assign layer_0[1311] = ~in[231] | (in[231] & in[120]); 
    assign layer_0[1312] = in[72]; 
    assign layer_0[1313] = ~(in[182] ^ in[150]); 
    assign layer_0[1314] = ~(in[90] ^ in[122]); 
    assign layer_0[1315] = ~in[22]; 
    assign layer_0[1316] = in[105] ^ in[125]; 
    assign layer_0[1317] = ~in[186] | (in[186] & in[70]); 
    assign layer_0[1318] = ~in[85] | (in[120] & in[85]); 
    assign layer_0[1319] = ~(in[196] ^ in[150]); 
    assign layer_0[1320] = ~(in[164] | in[182]); 
    assign layer_0[1321] = ~(in[204] | in[192]); 
    assign layer_0[1322] = in[194] ^ in[38]; 
    assign layer_0[1323] = ~(in[41] | in[99]); 
    assign layer_0[1324] = in[9]; 
    assign layer_0[1325] = ~in[121] | (in[121] & in[23]); 
    assign layer_0[1326] = ~(in[116] ^ in[118]); 
    assign layer_0[1327] = in[130] | in[115]; 
    assign layer_0[1328] = ~in[58] | (in[58] & in[181]); 
    assign layer_0[1329] = ~(in[101] ^ in[70]); 
    assign layer_0[1330] = ~(in[101] ^ in[99]); 
    assign layer_0[1331] = ~(in[228] | in[22]); 
    assign layer_0[1332] = ~(in[77] ^ in[45]); 
    assign layer_0[1333] = in[56] | in[228]; 
    assign layer_0[1334] = in[151] | in[166]; 
    assign layer_0[1335] = in[88] & ~in[43]; 
    assign layer_0[1336] = in[71] ^ in[36]; 
    assign layer_0[1337] = ~(in[236] | in[235]); 
    assign layer_0[1338] = in[183] | in[147]; 
    assign layer_0[1339] = ~(in[55] | in[72]); 
    assign layer_0[1340] = ~(in[188] ^ in[155]); 
    assign layer_0[1341] = ~(in[87] ^ in[56]); 
    assign layer_0[1342] = ~(in[105] ^ in[110]); 
    assign layer_0[1343] = in[206] ^ in[174]; 
    assign layer_0[1344] = in[24] ^ in[56]; 
    assign layer_0[1345] = in[133] & ~in[22]; 
    assign layer_0[1346] = ~(in[26] | in[196]); 
    assign layer_0[1347] = in[140] & ~in[75]; 
    assign layer_0[1348] = in[199] | in[54]; 
    assign layer_0[1349] = ~(in[61] ^ in[236]); 
    assign layer_0[1350] = ~(in[67] | in[83]); 
    assign layer_0[1351] = ~(in[160] | in[6]); 
    assign layer_0[1352] = ~in[103] | (in[220] & in[103]); 
    assign layer_0[1353] = in[130] ^ in[132]; 
    assign layer_0[1354] = in[90] | in[34]; 
    assign layer_0[1355] = ~in[215] | (in[247] & in[215]); 
    assign layer_0[1356] = in[165]; 
    assign layer_0[1357] = ~in[211]; 
    assign layer_0[1358] = in[70] ^ in[103]; 
    assign layer_0[1359] = in[56] & in[72]; 
    assign layer_0[1360] = ~(in[106] ^ in[153]); 
    assign layer_0[1361] = in[107] ^ in[121]; 
    assign layer_0[1362] = ~in[184]; 
    assign layer_0[1363] = in[198] ^ in[246]; 
    assign layer_0[1364] = ~(in[92] ^ in[53]); 
    assign layer_0[1365] = ~(in[173] | in[9]); 
    assign layer_0[1366] = ~in[53]; 
    assign layer_0[1367] = in[180] ^ in[182]; 
    assign layer_0[1368] = ~(in[29] | in[11]); 
    assign layer_0[1369] = ~in[170] | (in[249] & in[170]); 
    assign layer_0[1370] = in[218] ^ in[187]; 
    assign layer_0[1371] = in[169] ^ in[138]; 
    assign layer_0[1372] = in[171] ^ in[181]; 
    assign layer_0[1373] = in[196] ^ in[8]; 
    assign layer_0[1374] = ~(in[26] | in[25]); 
    assign layer_0[1375] = ~(in[129] ^ in[131]); 
    assign layer_0[1376] = in[205] | in[203]; 
    assign layer_0[1377] = ~(in[122] | in[156]); 
    assign layer_0[1378] = ~in[196]; 
    assign layer_0[1379] = in[39] ^ in[103]; 
    assign layer_0[1380] = ~(in[65] ^ in[34]); 
    assign layer_0[1381] = in[86] ^ in[100]; 
    assign layer_0[1382] = ~(in[24] | in[41]); 
    assign layer_0[1383] = ~(in[21] | in[137]); 
    assign layer_0[1384] = ~(in[163] | in[165]); 
    assign layer_0[1385] = in[150] ^ in[196]; 
    assign layer_0[1386] = in[54] ^ in[60]; 
    assign layer_0[1387] = ~(in[250] ^ in[248]); 
    assign layer_0[1388] = in[91] ^ in[93]; 
    assign layer_0[1389] = in[155] | in[124]; 
    assign layer_0[1390] = in[134] & in[153]; 
    assign layer_0[1391] = in[194] ^ in[196]; 
    assign layer_0[1392] = in[7] | in[163]; 
    assign layer_0[1393] = ~in[97]; 
    assign layer_0[1394] = ~in[76] | (in[106] & in[76]); 
    assign layer_0[1395] = in[117] ^ in[103]; 
    assign layer_0[1396] = ~(in[211] | in[233]); 
    assign layer_0[1397] = ~(in[24] ^ in[58]); 
    assign layer_0[1398] = ~in[105] | (in[68] & in[105]); 
    assign layer_0[1399] = in[59] & ~in[122]; 
    assign layer_0[1400] = ~in[117] | (in[117] & in[212]); 
    assign layer_0[1401] = ~(in[71] ^ in[85]); 
    assign layer_0[1402] = ~(in[102] ^ in[187]); 
    assign layer_0[1403] = in[66] ^ in[35]; 
    assign layer_0[1404] = in[164] | in[146]; 
    assign layer_0[1405] = in[120] & ~in[117]; 
    assign layer_0[1406] = ~(in[77] | in[234]); 
    assign layer_0[1407] = in[234] | in[245]; 
    assign layer_0[1408] = ~(in[59] ^ in[90]); 
    assign layer_0[1409] = in[157] | in[103]; 
    assign layer_0[1410] = ~(in[54] ^ in[199]); 
    assign layer_0[1411] = in[30] | in[110]; 
    assign layer_0[1412] = in[83]; 
    assign layer_0[1413] = in[230] ^ in[111]; 
    assign layer_0[1414] = in[232] & in[199]; 
    assign layer_0[1415] = ~in[182] | (in[182] & in[78]); 
    assign layer_0[1416] = in[170] & ~in[119]; 
    assign layer_0[1417] = in[202] & ~in[125]; 
    assign layer_0[1418] = ~(in[146] | in[145]); 
    assign layer_0[1419] = in[93] & ~in[120]; 
    assign layer_0[1420] = in[39] | in[87]; 
    assign layer_0[1421] = ~(in[186] | in[26]); 
    assign layer_0[1422] = ~in[77]; 
    assign layer_0[1423] = in[165] & ~in[248]; 
    assign layer_0[1424] = ~(in[119] | in[72]); 
    assign layer_0[1425] = in[99] ^ in[85]; 
    assign layer_0[1426] = in[198] ^ in[212]; 
    assign layer_0[1427] = in[106]; 
    assign layer_0[1428] = ~in[165] | (in[165] & in[172]); 
    assign layer_0[1429] = in[180] | in[178]; 
    assign layer_0[1430] = in[87] | in[105]; 
    assign layer_0[1431] = ~(in[221] | in[235]); 
    assign layer_0[1432] = in[244] | in[157]; 
    assign layer_0[1433] = ~(in[241] ^ in[151]); 
    assign layer_0[1434] = in[236] ^ in[205]; 
    assign layer_0[1435] = ~(in[218] | in[41]); 
    assign layer_0[1436] = ~(in[235] ^ in[186]); 
    assign layer_0[1437] = ~in[117]; 
    assign layer_0[1438] = in[88] ^ in[57]; 
    assign layer_0[1439] = in[74] ^ in[77]; 
    assign layer_0[1440] = in[231] & ~in[123]; 
    assign layer_0[1441] = ~(in[177] | in[8]); 
    assign layer_0[1442] = in[148]; 
    assign layer_0[1443] = ~(in[134] | in[149]); 
    assign layer_0[1444] = in[113] | in[123]; 
    assign layer_0[1445] = in[35] | in[218]; 
    assign layer_0[1446] = in[100] | in[85]; 
    assign layer_0[1447] = ~in[56] | (in[56] & in[198]); 
    assign layer_0[1448] = in[185] | in[140]; 
    assign layer_0[1449] = ~(in[136] ^ in[101]); 
    assign layer_0[1450] = in[174] | in[25]; 
    assign layer_0[1451] = in[104] & ~in[101]; 
    assign layer_0[1452] = in[70] ^ in[129]; 
    assign layer_0[1453] = ~(in[83] | in[53]); 
    assign layer_0[1454] = ~in[123] | (in[104] & in[123]); 
    assign layer_0[1455] = ~in[164]; 
    assign layer_0[1456] = in[76] ^ in[184]; 
    assign layer_0[1457] = ~(in[82] ^ in[178]); 
    assign layer_0[1458] = in[168] & ~in[139]; 
    assign layer_0[1459] = ~(in[89] ^ in[68]); 
    assign layer_0[1460] = in[57] & ~in[104]; 
    assign layer_0[1461] = in[100] & ~in[212]; 
    assign layer_0[1462] = ~in[72]; 
    assign layer_0[1463] = in[227] & ~in[251]; 
    assign layer_0[1464] = in[74] & ~in[100]; 
    assign layer_0[1465] = in[119] | in[163]; 
    assign layer_0[1466] = in[154]; 
    assign layer_0[1467] = ~(in[5] | in[92]); 
    assign layer_0[1468] = in[147]; 
    assign layer_0[1469] = ~(in[236] ^ in[8]); 
    assign layer_0[1470] = in[237] | in[169]; 
    assign layer_0[1471] = in[111] | in[109]; 
    assign layer_0[1472] = ~(in[117] | in[28]); 
    assign layer_0[1473] = in[119] | in[55]; 
    assign layer_0[1474] = ~in[8]; 
    assign layer_0[1475] = ~(in[52] ^ in[172]); 
    assign layer_0[1476] = in[150]; 
    assign layer_0[1477] = ~(in[183] ^ in[121]); 
    assign layer_0[1478] = in[83] ^ in[79]; 
    assign layer_0[1479] = in[40] ^ in[87]; 
    assign layer_0[1480] = in[185] | in[183]; 
    assign layer_0[1481] = in[189] | in[156]; 
    assign layer_0[1482] = ~(in[79] | in[47]); 
    assign layer_0[1483] = ~(in[108] ^ in[106]); 
    assign layer_0[1484] = ~in[217] | (in[217] & in[211]); 
    assign layer_0[1485] = ~(in[200] ^ in[196]); 
    assign layer_0[1486] = in[22] ^ in[136]; 
    assign layer_0[1487] = ~(in[40] ^ in[72]); 
    assign layer_0[1488] = in[202] ^ in[51]; 
    assign layer_0[1489] = in[58] | in[115]; 
    assign layer_0[1490] = in[71] ^ in[24]; 
    assign layer_0[1491] = in[213] | in[87]; 
    assign layer_0[1492] = in[250] ^ in[216]; 
    assign layer_0[1493] = in[101] & ~in[37]; 
    assign layer_0[1494] = in[147] ^ in[118]; 
    assign layer_0[1495] = in[103] ^ in[38]; 
    assign layer_0[1496] = in[39]; 
    assign layer_0[1497] = in[21] ^ in[162]; 
    assign layer_0[1498] = ~(in[253] | in[164]); 
    assign layer_0[1499] = in[145] | in[146]; 
    assign layer_0[1500] = ~(in[234] ^ in[187]); 
    assign layer_0[1501] = ~in[234] | (in[180] & in[234]); 
    assign layer_0[1502] = in[97] ^ in[73]; 
    assign layer_0[1503] = in[231] & ~in[152]; 
    assign layer_0[1504] = in[167] ^ in[100]; 
    assign layer_0[1505] = in[44] ^ in[62]; 
    assign layer_0[1506] = in[183] | in[164]; 
    assign layer_0[1507] = in[119] ^ in[166]; 
    assign layer_0[1508] = ~(in[165] ^ in[167]); 
    assign layer_0[1509] = in[170] ^ in[102]; 
    assign layer_0[1510] = in[180] & ~in[113]; 
    assign layer_0[1511] = ~(in[196] | in[216]); 
    assign layer_0[1512] = ~in[74] | (in[13] & in[74]); 
    assign layer_0[1513] = ~(in[40] ^ in[24]); 
    assign layer_0[1514] = in[22] ^ in[247]; 
    assign layer_0[1515] = ~in[168] | (in[168] & in[78]); 
    assign layer_0[1516] = in[73]; 
    assign layer_0[1517] = in[93] ^ in[66]; 
    assign layer_0[1518] = ~(in[200] ^ in[37]); 
    assign layer_0[1519] = in[73] ^ in[61]; 
    assign layer_0[1520] = in[66] ^ in[34]; 
    assign layer_0[1521] = ~(in[79] ^ in[30]); 
    assign layer_0[1522] = ~(in[135] ^ in[166]); 
    assign layer_0[1523] = in[73] & ~in[194]; 
    assign layer_0[1524] = ~in[133] | (in[133] & in[173]); 
    assign layer_0[1525] = in[129] ^ in[115]; 
    assign layer_0[1526] = ~(in[247] ^ in[250]); 
    assign layer_0[1527] = ~(in[247] ^ in[250]); 
    assign layer_0[1528] = in[165] ^ in[147]; 
    assign layer_0[1529] = in[98] | in[46]; 
    assign layer_0[1530] = ~in[75] | (in[29] & in[75]); 
    assign layer_0[1531] = in[63] ^ in[114]; 
    assign layer_0[1532] = in[23] ^ in[70]; 
    assign layer_0[1533] = in[173] ^ in[37]; 
    assign layer_0[1534] = ~in[56] | (in[60] & in[56]); 
    assign layer_0[1535] = in[152] & ~in[58]; 
    assign layer_0[1536] = in[106] ^ in[248]; 
    assign layer_0[1537] = in[247] ^ in[251]; 
    assign layer_0[1538] = in[120] & ~in[181]; 
    assign layer_0[1539] = in[69] ^ in[109]; 
    assign layer_0[1540] = in[231]; 
    assign layer_0[1541] = ~in[75] | (in[116] & in[75]); 
    assign layer_0[1542] = ~(in[107] ^ in[125]); 
    assign layer_0[1543] = in[99] & ~in[88]; 
    assign layer_0[1544] = in[229] ^ in[198]; 
    assign layer_0[1545] = in[147] & ~in[134]; 
    assign layer_0[1546] = in[82] | in[36]; 
    assign layer_0[1547] = in[152] & ~in[145]; 
    assign layer_0[1548] = in[54] & ~in[10]; 
    assign layer_0[1549] = in[195] ^ in[197]; 
    assign layer_0[1550] = in[11] & ~in[194]; 
    assign layer_0[1551] = in[109] ^ in[140]; 
    assign layer_0[1552] = ~(in[29] ^ in[63]); 
    assign layer_0[1553] = in[88]; 
    assign layer_0[1554] = in[179] | in[205]; 
    assign layer_0[1555] = ~(in[219] ^ in[235]); 
    assign layer_0[1556] = ~in[169]; 
    assign layer_0[1557] = in[104] ^ in[142]; 
    assign layer_0[1558] = ~in[244]; 
    assign layer_0[1559] = in[92] ^ in[95]; 
    assign layer_0[1560] = in[245] ^ in[251]; 
    assign layer_0[1561] = ~(in[170] ^ in[242]); 
    assign layer_0[1562] = ~(in[147] & in[130]); 
    assign layer_0[1563] = in[86] ^ in[41]; 
    assign layer_0[1564] = ~(in[117] ^ in[102]); 
    assign layer_0[1565] = in[164] ^ in[135]; 
    assign layer_0[1566] = in[142] ^ in[29]; 
    assign layer_0[1567] = in[210] ^ in[245]; 
    assign layer_0[1568] = ~in[120]; 
    assign layer_0[1569] = ~(in[108] ^ in[110]); 
    assign layer_0[1570] = ~(in[185] ^ in[167]); 
    assign layer_0[1571] = in[70] & ~in[212]; 
    assign layer_0[1572] = in[183] & ~in[176]; 
    assign layer_0[1573] = ~(in[124] | in[26]); 
    assign layer_0[1574] = in[182] & ~in[171]; 
    assign layer_0[1575] = in[121] & ~in[141]; 
    assign layer_0[1576] = in[115] ^ in[113]; 
    assign layer_0[1577] = ~in[7]; 
    assign layer_0[1578] = ~(in[150] ^ in[119]); 
    assign layer_0[1579] = in[53] | in[86]; 
    assign layer_0[1580] = ~(in[21] ^ in[53]); 
    assign layer_0[1581] = ~(in[202] | in[219]); 
    assign layer_0[1582] = ~(in[166] | in[163]); 
    assign layer_0[1583] = ~(in[184] | in[120]); 
    assign layer_0[1584] = ~(in[153] ^ in[218]); 
    assign layer_0[1585] = in[101] & ~in[22]; 
    assign layer_0[1586] = in[167] & ~in[156]; 
    assign layer_0[1587] = ~in[59] | (in[59] & in[243]); 
    assign layer_0[1588] = ~in[152] | (in[200] & in[152]); 
    assign layer_0[1589] = ~in[219] | (in[83] & in[219]); 
    assign layer_0[1590] = in[60] ^ in[45]; 
    assign layer_0[1591] = in[118] | in[131]; 
    assign layer_0[1592] = ~(in[85] ^ in[52]); 
    assign layer_0[1593] = ~(in[176] | in[137]); 
    assign layer_0[1594] = in[177] | in[99]; 
    assign layer_0[1595] = in[76] | in[75]; 
    assign layer_0[1596] = ~(in[8] | in[22]); 
    assign layer_0[1597] = ~(in[232] & in[184]); 
    assign layer_0[1598] = in[164] ^ in[182]; 
    assign layer_0[1599] = ~in[198] | (in[198] & in[92]); 
    // Layer 1 ============================================================
    assign out[0] = ~(layer_0[1587] ^ layer_0[830]); 
    assign out[1] = ~(layer_0[82] ^ layer_0[1240]); 
    assign out[2] = ~(layer_0[916] ^ layer_0[715]); 
    assign out[3] = layer_0[968]; 
    assign out[4] = ~(layer_0[464] ^ layer_0[1017]); 
    assign out[5] = layer_0[417] & layer_0[569]; 
    assign out[6] = layer_0[650] & ~layer_0[1111]; 
    assign out[7] = ~(layer_0[1234] ^ layer_0[1572]); 
    assign out[8] = layer_0[614] & ~layer_0[524]; 
    assign out[9] = layer_0[54] | layer_0[416]; 
    assign out[10] = layer_0[572] & ~layer_0[24]; 
    assign out[11] = layer_0[301] & ~layer_0[426]; 
    assign out[12] = ~(layer_0[622] & layer_0[100]); 
    assign out[13] = ~layer_0[865]; 
    assign out[14] = layer_0[378]; 
    assign out[15] = ~layer_0[1304]; 
    assign out[16] = ~layer_0[37]; 
    assign out[17] = ~(layer_0[194] ^ layer_0[1570]); 
    assign out[18] = layer_0[940] & ~layer_0[1418]; 
    assign out[19] = ~layer_0[190]; 
    assign out[20] = ~layer_0[1016]; 
    assign out[21] = layer_0[245] & ~layer_0[926]; 
    assign out[22] = ~(layer_0[654] & layer_0[911]); 
    assign out[23] = ~layer_0[1255] | (layer_0[1495] & layer_0[1255]); 
    assign out[24] = ~layer_0[649]; 
    assign out[25] = layer_0[276] & layer_0[211]; 
    assign out[26] = layer_0[998] & layer_0[10]; 
    assign out[27] = ~layer_0[246]; 
    assign out[28] = layer_0[898] & layer_0[651]; 
    assign out[29] = layer_0[1085] | layer_0[73]; 
    assign out[30] = layer_0[481] | layer_0[828]; 
    assign out[31] = layer_0[103] & ~layer_0[1330]; 
    assign out[32] = ~layer_0[886]; 
    assign out[33] = layer_0[534] & ~layer_0[783]; 
    assign out[34] = layer_0[1568] & ~layer_0[1560]; 
    assign out[35] = ~layer_0[324]; 
    assign out[36] = layer_0[327] ^ layer_0[226]; 
    assign out[37] = layer_0[338] ^ layer_0[613]; 
    assign out[38] = ~layer_0[1060]; 
    assign out[39] = ~layer_0[1273]; 
    assign out[40] = layer_0[75] & ~layer_0[396]; 
    assign out[41] = ~layer_0[1569]; 
    assign out[42] = ~(layer_0[158] ^ layer_0[763]); 
    assign out[43] = layer_0[733] ^ layer_0[133]; 
    assign out[44] = layer_0[1522] & ~layer_0[733]; 
    assign out[45] = ~layer_0[838]; 
    assign out[46] = ~layer_0[1378] | (layer_0[1378] & layer_0[1305]); 
    assign out[47] = ~layer_0[444]; 
    assign out[48] = layer_0[677] & ~layer_0[627]; 
    assign out[49] = ~layer_0[679]; 
    assign out[50] = layer_0[1185] & layer_0[213]; 
    assign out[51] = ~layer_0[743]; 
    assign out[52] = layer_0[821]; 
    assign out[53] = ~layer_0[163] | (layer_0[748] & layer_0[163]); 
    assign out[54] = layer_0[1063]; 
    assign out[55] = ~layer_0[413]; 
    assign out[56] = layer_0[1509] ^ layer_0[374]; 
    assign out[57] = layer_0[384] & ~layer_0[815]; 
    assign out[58] = layer_0[319] & ~layer_0[1159]; 
    assign out[59] = ~layer_0[861]; 
    assign out[60] = ~(layer_0[244] ^ layer_0[1558]); 
    assign out[61] = ~(layer_0[1283] & layer_0[715]); 
    assign out[62] = ~(layer_0[450] | layer_0[387]); 
    assign out[63] = layer_0[1503] ^ layer_0[381]; 
    assign out[64] = layer_0[1314]; 
    assign out[65] = layer_0[1257] ^ layer_0[248]; 
    assign out[66] = layer_0[1327] ^ layer_0[924]; 
    assign out[67] = layer_0[1383] & layer_0[1500]; 
    assign out[68] = ~layer_0[1369] | (layer_0[1369] & layer_0[1165]); 
    assign out[69] = layer_0[1152] & layer_0[689]; 
    assign out[70] = ~layer_0[950]; 
    assign out[71] = layer_0[475]; 
    assign out[72] = ~(layer_0[801] ^ layer_0[943]); 
    assign out[73] = ~layer_0[1486]; 
    assign out[74] = ~layer_0[794] | (layer_0[1583] & layer_0[794]); 
    assign out[75] = layer_0[1578]; 
    assign out[76] = ~(layer_0[1065] ^ layer_0[984]); 
    assign out[77] = layer_0[40]; 
    assign out[78] = ~layer_0[11] | (layer_0[11] & layer_0[358]); 
    assign out[79] = ~(layer_0[267] ^ layer_0[1088]); 
    assign out[80] = ~(layer_0[981] ^ layer_0[1046]); 
    assign out[81] = ~(layer_0[1438] ^ layer_0[1120]); 
    assign out[82] = layer_0[4]; 
    assign out[83] = ~(layer_0[1172] ^ layer_0[227]); 
    assign out[84] = layer_0[900] & layer_0[1057]; 
    assign out[85] = layer_0[980]; 
    assign out[86] = ~(layer_0[551] | layer_0[1023]); 
    assign out[87] = layer_0[456] & layer_0[9]; 
    assign out[88] = ~(layer_0[139] ^ layer_0[1068]); 
    assign out[89] = layer_0[101] & layer_0[985]; 
    assign out[90] = layer_0[1205] ^ layer_0[253]; 
    assign out[91] = ~(layer_0[938] ^ layer_0[235]); 
    assign out[92] = ~layer_0[1197]; 
    assign out[93] = layer_0[171] ^ layer_0[1039]; 
    assign out[94] = layer_0[796]; 
    assign out[95] = layer_0[1491] & ~layer_0[655]; 
    assign out[96] = ~(layer_0[1311] | layer_0[541]); 
    assign out[97] = layer_0[302] & ~layer_0[1371]; 
    assign out[98] = ~(layer_0[212] & layer_0[854]); 
    assign out[99] = layer_0[442]; 
    assign out[100] = layer_0[117] & ~layer_0[1547]; 
    assign out[101] = ~(layer_0[698] | layer_0[359]); 
    assign out[102] = layer_0[469]; 
    assign out[103] = ~layer_0[1092] | (layer_0[548] & layer_0[1092]); 
    assign out[104] = layer_0[1203] & ~layer_0[636]; 
    assign out[105] = layer_0[1426]; 
    assign out[106] = ~(layer_0[563] ^ layer_0[947]); 
    assign out[107] = ~(layer_0[364] ^ layer_0[1430]); 
    assign out[108] = layer_0[168] & ~layer_0[597]; 
    assign out[109] = layer_0[1593] & ~layer_0[630]; 
    assign out[110] = layer_0[177]; 
    assign out[111] = layer_0[485] ^ layer_0[1432]; 
    assign out[112] = ~(layer_0[54] ^ layer_0[805]); 
    assign out[113] = ~(layer_0[1399] ^ layer_0[1318]); 
    assign out[114] = ~(layer_0[96] & layer_0[910]); 
    assign out[115] = layer_0[729] & ~layer_0[69]; 
    assign out[116] = layer_0[1383] & layer_0[680]; 
    assign out[117] = ~layer_0[364]; 
    assign out[118] = ~layer_0[745] | (layer_0[781] & layer_0[745]); 
    assign out[119] = layer_0[192] ^ layer_0[500]; 
    assign out[120] = layer_0[672]; 
    assign out[121] = layer_0[62] | layer_0[775]; 
    assign out[122] = layer_0[311] & ~layer_0[584]; 
    assign out[123] = layer_0[1419] | layer_0[170]; 
    assign out[124] = layer_0[1489] & ~layer_0[874]; 
    assign out[125] = ~(layer_0[758] ^ layer_0[1027]); 
    assign out[126] = layer_0[1362] ^ layer_0[1007]; 
    assign out[127] = ~(layer_0[810] ^ layer_0[118]); 
    assign out[128] = layer_0[1534] ^ layer_0[1067]; 
    assign out[129] = layer_0[711] ^ layer_0[156]; 
    assign out[130] = ~(layer_0[1181] ^ layer_0[1414]); 
    assign out[131] = layer_0[452] & ~layer_0[14]; 
    assign out[132] = layer_0[1031] & ~layer_0[187]; 
    assign out[133] = ~(layer_0[983] | layer_0[281]); 
    assign out[134] = layer_0[1530] & ~layer_0[65]; 
    assign out[135] = ~layer_0[423] | (layer_0[108] & layer_0[423]); 
    assign out[136] = ~(layer_0[179] ^ layer_0[660]); 
    assign out[137] = layer_0[184]; 
    assign out[138] = layer_0[765] ^ layer_0[195]; 
    assign out[139] = layer_0[1439] ^ layer_0[467]; 
    assign out[140] = ~layer_0[495]; 
    assign out[141] = ~(layer_0[760] ^ layer_0[17]); 
    assign out[142] = ~(layer_0[127] ^ layer_0[395]); 
    assign out[143] = layer_0[568]; 
    assign out[144] = ~(layer_0[503] ^ layer_0[1420]); 
    assign out[145] = layer_0[707] ^ layer_0[1384]; 
    assign out[146] = layer_0[1553] ^ layer_0[575]; 
    assign out[147] = ~(layer_0[1033] ^ layer_0[1124]); 
    assign out[148] = layer_0[554] & layer_0[120]; 
    assign out[149] = layer_0[373] & layer_0[232]; 
    assign out[150] = layer_0[525] & ~layer_0[1217]; 
    assign out[151] = layer_0[1180] & ~layer_0[330]; 
    assign out[152] = layer_0[601]; 
    assign out[153] = layer_0[1014] & ~layer_0[1449]; 
    assign out[154] = layer_0[1182] & ~layer_0[791]; 
    assign out[155] = layer_0[1491] & layer_0[661]; 
    assign out[156] = ~(layer_0[1129] ^ layer_0[785]); 
    assign out[157] = layer_0[862] & ~layer_0[859]; 
    assign out[158] = layer_0[1484] & ~layer_0[134]; 
    assign out[159] = ~(layer_0[234] ^ layer_0[351]); 
    assign out[160] = ~(layer_0[785] ^ layer_0[708]); 
    assign out[161] = layer_0[1137] ^ layer_0[1431]; 
    assign out[162] = layer_0[94] & layer_0[1580]; 
    assign out[163] = ~(layer_0[992] | layer_0[953]); 
    assign out[164] = ~(layer_0[948] ^ layer_0[993]); 
    assign out[165] = layer_0[19] ^ layer_0[1266]; 
    assign out[166] = layer_0[1317] & ~layer_0[1532]; 
    assign out[167] = layer_0[440] ^ layer_0[729]; 
    assign out[168] = layer_0[1265] & ~layer_0[18]; 
    assign out[169] = layer_0[689] & ~layer_0[1459]; 
    assign out[170] = ~(layer_0[184] ^ layer_0[1467]); 
    assign out[171] = ~(layer_0[804] | layer_0[1597]); 
    assign out[172] = ~(layer_0[40] | layer_0[1075]); 
    assign out[173] = layer_0[601] | layer_0[915]; 
    assign out[174] = layer_0[1091] & layer_0[1105]; 
    assign out[175] = ~layer_0[332] | (layer_0[131] & layer_0[332]); 
    assign out[176] = layer_0[1463] ^ layer_0[482]; 
    assign out[177] = ~layer_0[354]; 
    assign out[178] = ~(layer_0[1594] | layer_0[209]); 
    assign out[179] = layer_0[838] & layer_0[1422]; 
    assign out[180] = ~(layer_0[137] ^ layer_0[614]); 
    assign out[181] = layer_0[912] ^ layer_0[923]; 
    assign out[182] = ~(layer_0[1389] | layer_0[857]); 
    assign out[183] = layer_0[23] & ~layer_0[1478]; 
    assign out[184] = layer_0[419] & layer_0[1117]; 
    assign out[185] = ~(layer_0[134] ^ layer_0[948]); 
    assign out[186] = layer_0[994] & ~layer_0[722]; 
    assign out[187] = ~(layer_0[242] ^ layer_0[723]); 
    assign out[188] = layer_0[1006] & ~layer_0[1288]; 
    assign out[189] = layer_0[323]; 
    assign out[190] = ~layer_0[88]; 
    assign out[191] = layer_0[458] & layer_0[1035]; 
    assign out[192] = layer_0[1577] ^ layer_0[996]; 
    assign out[193] = layer_0[231] ^ layer_0[98]; 
    assign out[194] = layer_0[108] & ~layer_0[288]; 
    assign out[195] = ~layer_0[593]; 
    assign out[196] = layer_0[1287] | layer_0[1550]; 
    assign out[197] = layer_0[606] ^ layer_0[183]; 
    assign out[198] = layer_0[224] ^ layer_0[1529]; 
    assign out[199] = layer_0[439]; 
    assign out[200] = ~(layer_0[410] | layer_0[1322]); 
    assign out[201] = layer_0[780]; 
    assign out[202] = layer_0[337] & ~layer_0[811]; 
    assign out[203] = layer_0[1223] | layer_0[517]; 
    assign out[204] = ~(layer_0[1529] ^ layer_0[206]); 
    assign out[205] = layer_0[25] ^ layer_0[1022]; 
    assign out[206] = ~layer_0[398]; 
    assign out[207] = layer_0[1515] ^ layer_0[833]; 
    assign out[208] = layer_0[687] ^ layer_0[401]; 
    assign out[209] = layer_0[1509] ^ layer_0[79]; 
    assign out[210] = ~(layer_0[1205] | layer_0[593]); 
    assign out[211] = ~layer_0[155]; 
    assign out[212] = layer_0[453] | layer_0[1218]; 
    assign out[213] = ~(layer_0[744] ^ layer_0[1054]); 
    assign out[214] = layer_0[1073]; 
    assign out[215] = layer_0[197]; 
    assign out[216] = ~(layer_0[95] | layer_0[1045]); 
    assign out[217] = ~(layer_0[888] ^ layer_0[1369]); 
    assign out[218] = ~(layer_0[1325] ^ layer_0[179]); 
    assign out[219] = ~(layer_0[1551] | layer_0[1368]); 
    assign out[220] = layer_0[1292] & ~layer_0[727]; 
    assign out[221] = ~layer_0[300]; 
    assign out[222] = ~(layer_0[1485] ^ layer_0[1546]); 
    assign out[223] = layer_0[628] ^ layer_0[206]; 
    assign out[224] = layer_0[764] ^ layer_0[326]; 
    assign out[225] = layer_0[1124] ^ layer_0[411]; 
    assign out[226] = ~(layer_0[1201] ^ layer_0[545]); 
    assign out[227] = ~layer_0[243]; 
    assign out[228] = layer_0[1022] & ~layer_0[139]; 
    assign out[229] = layer_0[362]; 
    assign out[230] = layer_0[521] & ~layer_0[339]; 
    assign out[231] = layer_0[487] | layer_0[1451]; 
    assign out[232] = layer_0[600]; 
    assign out[233] = layer_0[995] & layer_0[194]; 
    assign out[234] = ~(layer_0[834] ^ layer_0[314]); 
    assign out[235] = layer_0[106] | layer_0[1434]; 
    assign out[236] = layer_0[1188] & ~layer_0[764]; 
    assign out[237] = ~layer_0[1101]; 
    assign out[238] = layer_0[884]; 
    assign out[239] = layer_0[1094] ^ layer_0[1535]; 
    assign out[240] = layer_0[1102] & layer_0[960]; 
    assign out[241] = layer_0[1284] & ~layer_0[666]; 
    assign out[242] = ~(layer_0[1297] & layer_0[1555]); 
    assign out[243] = layer_0[222] & ~layer_0[1025]; 
    assign out[244] = layer_0[1024]; 
    assign out[245] = ~layer_0[1215] | (layer_0[1215] & layer_0[578]); 
    assign out[246] = layer_0[445] & ~layer_0[611]; 
    assign out[247] = ~layer_0[1153]; 
    assign out[248] = ~(layer_0[1034] ^ layer_0[1372]); 
    assign out[249] = layer_0[1232] ^ layer_0[110]; 
    assign out[250] = ~(layer_0[688] ^ layer_0[1082]); 
    assign out[251] = layer_0[803] & layer_0[422]; 
    assign out[252] = layer_0[265] ^ layer_0[975]; 
    assign out[253] = layer_0[507] ^ layer_0[1118]; 
    assign out[254] = layer_0[887] ^ layer_0[1015]; 
    assign out[255] = ~layer_0[1175]; 
    assign out[256] = layer_0[674]; 
    assign out[257] = ~layer_0[590] | (layer_0[902] & layer_0[590]); 
    assign out[258] = layer_0[589]; 
    assign out[259] = ~layer_0[160] | (layer_0[3] & layer_0[160]); 
    assign out[260] = ~(layer_0[880] | layer_0[1381]); 
    assign out[261] = ~(layer_0[1511] & layer_0[1407]); 
    assign out[262] = ~layer_0[1276]; 
    assign out[263] = layer_0[582]; 
    assign out[264] = layer_0[1326] & layer_0[1215]; 
    assign out[265] = ~layer_0[1156] | (layer_0[1329] & layer_0[1156]); 
    assign out[266] = ~(layer_0[112] ^ layer_0[1575]); 
    assign out[267] = ~layer_0[799] | (layer_0[932] & layer_0[799]); 
    assign out[268] = layer_0[1330] & ~layer_0[377]; 
    assign out[269] = layer_0[315]; 
    assign out[270] = ~layer_0[741] | (layer_0[741] & layer_0[1497]); 
    assign out[271] = layer_0[461] & ~layer_0[1537]; 
    assign out[272] = ~layer_0[1565]; 
    assign out[273] = layer_0[1545] ^ layer_0[1048]; 
    assign out[274] = ~layer_0[1531]; 
    assign out[275] = ~(layer_0[651] & layer_0[648]); 
    assign out[276] = ~layer_0[175] | (layer_0[585] & layer_0[175]); 
    assign out[277] = layer_0[1047] & ~layer_0[573]; 
    assign out[278] = layer_0[410] & ~layer_0[22]; 
    assign out[279] = layer_0[1003] & layer_0[445]; 
    assign out[280] = ~layer_0[205]; 
    assign out[281] = ~layer_0[86]; 
    assign out[282] = layer_0[58] | layer_0[240]; 
    assign out[283] = ~(layer_0[109] & layer_0[1214]); 
    assign out[284] = layer_0[1114] ^ layer_0[242]; 
    assign out[285] = layer_0[813] ^ layer_0[1092]; 
    assign out[286] = ~(layer_0[305] & layer_0[205]); 
    assign out[287] = ~layer_0[1500]; 
    assign out[288] = layer_0[64]; 
    assign out[289] = layer_0[1462] ^ layer_0[1374]; 
    assign out[290] = ~layer_0[983]; 
    assign out[291] = layer_0[800] & layer_0[1051]; 
    assign out[292] = ~layer_0[1040]; 
    assign out[293] = ~(layer_0[165] ^ layer_0[556]); 
    assign out[294] = layer_0[1074]; 
    assign out[295] = ~(layer_0[793] ^ layer_0[284]); 
    assign out[296] = ~(layer_0[1260] & layer_0[653]); 
    assign out[297] = layer_0[608]; 
    assign out[298] = ~(layer_0[844] ^ layer_0[628]); 
    assign out[299] = layer_0[539] & layer_0[484]; 
    assign out[300] = ~(layer_0[1142] ^ layer_0[605]); 
    assign out[301] = layer_0[1456]; 
    assign out[302] = ~(layer_0[477] ^ layer_0[185]); 
    assign out[303] = layer_0[1528] & layer_0[571]; 
    assign out[304] = layer_0[649]; 
    assign out[305] = ~(layer_0[326] & layer_0[1030]); 
    assign out[306] = layer_0[1158] & ~layer_0[483]; 
    assign out[307] = layer_0[1192] ^ layer_0[1155]; 
    assign out[308] = layer_0[1589] ^ layer_0[744]; 
    assign out[309] = ~layer_0[1011] | (layer_0[906] & layer_0[1011]); 
    assign out[310] = layer_0[1191] ^ layer_0[370]; 
    assign out[311] = layer_0[522] ^ layer_0[1352]; 
    assign out[312] = layer_0[1343] & ~layer_0[566]; 
    assign out[313] = layer_0[865]; 
    assign out[314] = ~layer_0[1143] | (layer_0[1143] & layer_0[133]); 
    assign out[315] = layer_0[1370]; 
    assign out[316] = ~layer_0[1557]; 
    assign out[317] = layer_0[407] & layer_0[1230]; 
    assign out[318] = ~(layer_0[847] ^ layer_0[295]); 
    assign out[319] = ~layer_0[111]; 
    assign out[320] = ~(layer_0[49] & layer_0[1551]); 
    assign out[321] = layer_0[27]; 
    assign out[322] = ~layer_0[1584]; 
    assign out[323] = ~(layer_0[225] ^ layer_0[1596]); 
    assign out[324] = layer_0[512]; 
    assign out[325] = ~layer_0[1525]; 
    assign out[326] = layer_0[1402] & layer_0[1025]; 
    assign out[327] = ~(layer_0[573] ^ layer_0[945]); 
    assign out[328] = ~(layer_0[49] & layer_0[430]); 
    assign out[329] = layer_0[817] | layer_0[1434]; 
    assign out[330] = layer_0[979] ^ layer_0[1411]; 
    assign out[331] = ~(layer_0[41] ^ layer_0[188]); 
    assign out[332] = layer_0[1599] ^ layer_0[367]; 
    assign out[333] = layer_0[1441] ^ layer_0[882]; 
    assign out[334] = layer_0[1269] | layer_0[712]; 
    assign out[335] = ~(layer_0[1274] & layer_0[702]); 
    assign out[336] = layer_0[1302] ^ layer_0[84]; 
    assign out[337] = layer_0[18] ^ layer_0[35]; 
    assign out[338] = layer_0[180] & layer_0[294]; 
    assign out[339] = ~(layer_0[647] ^ layer_0[448]); 
    assign out[340] = layer_0[114] ^ layer_0[918]; 
    assign out[341] = ~(layer_0[428] & layer_0[1285]); 
    assign out[342] = layer_0[1314]; 
    assign out[343] = ~layer_0[431] | (layer_0[713] & layer_0[431]); 
    assign out[344] = layer_0[1558] & ~layer_0[7]; 
    assign out[345] = ~(layer_0[774] ^ layer_0[353]); 
    assign out[346] = ~layer_0[669] | (layer_0[655] & layer_0[669]); 
    assign out[347] = ~layer_0[129] | (layer_0[129] & layer_0[1397]); 
    assign out[348] = ~(layer_0[196] & layer_0[1351]); 
    assign out[349] = layer_0[1209] ^ layer_0[73]; 
    assign out[350] = layer_0[1145] & layer_0[1326]; 
    assign out[351] = ~(layer_0[978] ^ layer_0[747]); 
    assign out[352] = layer_0[1406] | layer_0[61]; 
    assign out[353] = ~layer_0[1175] | (layer_0[1175] & layer_0[810]); 
    assign out[354] = layer_0[693]; 
    assign out[355] = layer_0[373]; 
    assign out[356] = layer_0[959] & ~layer_0[483]; 
    assign out[357] = layer_0[602] ^ layer_0[1258]; 
    assign out[358] = layer_0[1019] ^ layer_0[1058]; 
    assign out[359] = layer_0[727]; 
    assign out[360] = ~(layer_0[1395] ^ layer_0[1499]); 
    assign out[361] = layer_0[1003] & ~layer_0[1049]; 
    assign out[362] = layer_0[398]; 
    assign out[363] = ~(layer_0[1023] ^ layer_0[69]); 
    assign out[364] = ~(layer_0[1089] ^ layer_0[565]); 
    assign out[365] = ~(layer_0[848] ^ layer_0[1405]); 
    assign out[366] = ~layer_0[1457] | (layer_0[1549] & layer_0[1457]); 
    assign out[367] = ~(layer_0[501] | layer_0[1421]); 
    assign out[368] = ~(layer_0[1446] ^ layer_0[623]); 
    assign out[369] = ~layer_0[404]; 
    assign out[370] = ~(layer_0[702] ^ layer_0[893]); 
    assign out[371] = layer_0[250] | layer_0[58]; 
    assign out[372] = layer_0[429] | layer_0[141]; 
    assign out[373] = ~(layer_0[8] ^ layer_0[1204]); 
    assign out[374] = layer_0[1189] & ~layer_0[385]; 
    assign out[375] = layer_0[1056] & layer_0[1526]; 
    assign out[376] = ~layer_0[1289] | (layer_0[1289] & layer_0[1423]); 
    assign out[377] = layer_0[1398]; 
    assign out[378] = ~(layer_0[33] | layer_0[1538]); 
    assign out[379] = layer_0[999] & layer_0[1332]; 
    assign out[380] = layer_0[388]; 
    assign out[381] = ~layer_0[1286] | (layer_0[1286] & layer_0[496]); 
    assign out[382] = layer_0[820]; 
    assign out[383] = layer_0[1363]; 
    assign out[384] = layer_0[1182]; 
    assign out[385] = layer_0[420] & layer_0[57]; 
    assign out[386] = layer_0[788]; 
    assign out[387] = layer_0[741] & ~layer_0[432]; 
    assign out[388] = layer_0[1127] & ~layer_0[1449]; 
    assign out[389] = ~layer_0[1319]; 
    assign out[390] = layer_0[915] ^ layer_0[1417]; 
    assign out[391] = layer_0[494]; 
    assign out[392] = ~layer_0[987] | (layer_0[425] & layer_0[987]); 
    assign out[393] = layer_0[622]; 
    assign out[394] = layer_0[835]; 
    assign out[395] = layer_0[1226]; 
    assign out[396] = layer_0[474] & ~layer_0[1176]; 
    assign out[397] = ~layer_0[626]; 
    assign out[398] = ~layer_0[754] | (layer_0[1144] & layer_0[754]); 
    assign out[399] = layer_0[141]; 
    assign out[400] = layer_0[1262] & layer_0[555]; 
    assign out[401] = layer_0[1282]; 
    assign out[402] = ~(layer_0[872] ^ layer_0[37]); 
    assign out[403] = layer_0[56] ^ layer_0[697]; 
    assign out[404] = ~layer_0[1416]; 
    assign out[405] = ~(layer_0[956] & layer_0[672]); 
    assign out[406] = layer_0[309] ^ layer_0[1110]; 
    assign out[407] = layer_0[1349] ^ layer_0[967]; 
    assign out[408] = layer_0[603] & ~layer_0[332]; 
    assign out[409] = ~layer_0[1159]; 
    assign out[410] = layer_0[751] & ~layer_0[1061]; 
    assign out[411] = layer_0[486]; 
    assign out[412] = layer_0[877] & ~layer_0[385]; 
    assign out[413] = ~(layer_0[812] ^ layer_0[901]); 
    assign out[414] = ~(layer_0[1572] & layer_0[1380]); 
    assign out[415] = layer_0[819] & ~layer_0[557]; 
    assign out[416] = ~layer_0[1351]; 
    assign out[417] = layer_0[140] & ~layer_0[1079]; 
    assign out[418] = layer_0[888] ^ layer_0[84]; 
    assign out[419] = ~layer_0[1264]; 
    assign out[420] = layer_0[1187] ^ layer_0[503]; 
    assign out[421] = layer_0[964]; 
    assign out[422] = layer_0[1280] ^ layer_0[360]; 
    assign out[423] = layer_0[629]; 
    assign out[424] = layer_0[610]; 
    assign out[425] = ~(layer_0[876] | layer_0[2]); 
    assign out[426] = ~(layer_0[971] | layer_0[29]); 
    assign out[427] = layer_0[531] | layer_0[1519]; 
    assign out[428] = layer_0[972] | layer_0[1536]; 
    assign out[429] = ~(layer_0[505] & layer_0[488]); 
    assign out[430] = layer_0[788] & ~layer_0[1140]; 
    assign out[431] = ~(layer_0[1354] ^ layer_0[826]); 
    assign out[432] = ~(layer_0[379] ^ layer_0[1195]); 
    assign out[433] = layer_0[367] ^ layer_0[771]; 
    assign out[434] = layer_0[150] ^ layer_0[374]; 
    assign out[435] = layer_0[157] & ~layer_0[1235]; 
    assign out[436] = ~(layer_0[1139] ^ layer_0[814]); 
    assign out[437] = ~(layer_0[1327] ^ layer_0[1585]); 
    assign out[438] = ~(layer_0[93] ^ layer_0[1128]); 
    assign out[439] = layer_0[291] & ~layer_0[67]; 
    assign out[440] = layer_0[671]; 
    assign out[441] = ~(layer_0[665] | layer_0[1381]); 
    assign out[442] = layer_0[552] & ~layer_0[876]; 
    assign out[443] = layer_0[889]; 
    assign out[444] = ~layer_0[1336]; 
    assign out[445] = layer_0[1248] | layer_0[1147]; 
    assign out[446] = ~(layer_0[455] ^ layer_0[901]); 
    assign out[447] = ~(layer_0[10] ^ layer_0[912]); 
    assign out[448] = ~(layer_0[1050] | layer_0[1412]); 
    assign out[449] = ~(layer_0[424] ^ layer_0[1220]); 
    assign out[450] = layer_0[1394]; 
    assign out[451] = layer_0[721] & layer_0[15]; 
    assign out[452] = ~layer_0[274]; 
    assign out[453] = layer_0[1245]; 
    assign out[454] = layer_0[1321] ^ layer_0[1474]; 
    assign out[455] = layer_0[1305] ^ layer_0[145]; 
    assign out[456] = layer_0[260] & ~layer_0[1069]; 
    assign out[457] = ~layer_0[871]; 
    assign out[458] = ~layer_0[806]; 
    assign out[459] = ~(layer_0[609] ^ layer_0[380]); 
    assign out[460] = ~(layer_0[1279] ^ layer_0[360]); 
    assign out[461] = ~layer_0[739]; 
    assign out[462] = ~(layer_0[1530] | layer_0[328]); 
    assign out[463] = ~(layer_0[1219] ^ layer_0[1588]); 
    assign out[464] = layer_0[85] & layer_0[646]; 
    assign out[465] = ~(layer_0[583] ^ layer_0[1299]); 
    assign out[466] = ~layer_0[1128] | (layer_0[1516] & layer_0[1128]); 
    assign out[467] = layer_0[1005] & ~layer_0[841]; 
    assign out[468] = ~layer_0[1240]; 
    assign out[469] = ~layer_0[1291] | (layer_0[1291] & layer_0[612]); 
    assign out[470] = ~(layer_0[236] ^ layer_0[595]); 
    assign out[471] = layer_0[718] ^ layer_0[1306]; 
    assign out[472] = layer_0[1492]; 
    assign out[473] = layer_0[19] ^ layer_0[9]; 
    assign out[474] = layer_0[1040] & ~layer_0[1425]; 
    assign out[475] = layer_0[873] ^ layer_0[1437]; 
    assign out[476] = layer_0[574] & layer_0[52]; 
    assign out[477] = ~(layer_0[154] ^ layer_0[942]); 
    assign out[478] = layer_0[1520]; 
    assign out[479] = ~layer_0[144]; 
    assign out[480] = ~layer_0[1518]; 
    assign out[481] = ~(layer_0[1206] ^ layer_0[631]); 
    assign out[482] = layer_0[855] | layer_0[173]; 
    assign out[483] = layer_0[65] ^ layer_0[307]; 
    assign out[484] = layer_0[594] ^ layer_0[678]; 
    assign out[485] = ~(layer_0[963] ^ layer_0[1160]); 
    assign out[486] = ~layer_0[1442] | (layer_0[1442] & layer_0[746]); 
    assign out[487] = layer_0[1401] & ~layer_0[204]; 
    assign out[488] = layer_0[261] & layer_0[551]; 
    assign out[489] = layer_0[779] ^ layer_0[1134]; 
    assign out[490] = layer_0[759] ^ layer_0[520]; 
    assign out[491] = layer_0[119] & ~layer_0[319]; 
    assign out[492] = layer_0[1007]; 
    assign out[493] = layer_0[762] & ~layer_0[832]; 
    assign out[494] = ~(layer_0[1014] | layer_0[240]); 
    assign out[495] = layer_0[600] ^ layer_0[1237]; 
    assign out[496] = layer_0[120]; 
    assign out[497] = layer_0[571] & ~layer_0[21]; 
    assign out[498] = ~(layer_0[1581] | layer_0[1029]); 
    assign out[499] = layer_0[618] & layer_0[855]; 
    assign out[500] = layer_0[1077]; 
    assign out[501] = layer_0[265]; 
    assign out[502] = ~(layer_0[1044] ^ layer_0[633]); 
    assign out[503] = ~(layer_0[1076] | layer_0[1339]); 
    assign out[504] = layer_0[1365] ^ layer_0[372]; 
    assign out[505] = layer_0[1016] ^ layer_0[449]; 
    assign out[506] = layer_0[43] & ~layer_0[973]; 
    assign out[507] = ~(layer_0[1380] & layer_0[951]); 
    assign out[508] = ~layer_0[1490]; 
    assign out[509] = layer_0[1239] & ~layer_0[341]; 
    assign out[510] = layer_0[761] ^ layer_0[502]; 
    assign out[511] = ~layer_0[1227]; 
    assign out[512] = ~layer_0[693]; 
    assign out[513] = layer_0[340] & ~layer_0[1539]; 
    assign out[514] = layer_0[1037]; 
    assign out[515] = layer_0[585]; 
    assign out[516] = layer_0[264] ^ layer_0[321]; 
    assign out[517] = layer_0[1171] ^ layer_0[767]; 
    assign out[518] = layer_0[952] & ~layer_0[795]; 
    assign out[519] = ~layer_0[647] | (layer_0[647] & layer_0[708]); 
    assign out[520] = ~(layer_0[318] & layer_0[480]); 
    assign out[521] = ~(layer_0[104] ^ layer_0[204]); 
    assign out[522] = ~(layer_0[437] ^ layer_0[1039]); 
    assign out[523] = layer_0[138] | layer_0[1543]; 
    assign out[524] = ~(layer_0[1401] & layer_0[1127]); 
    assign out[525] = ~layer_0[400]; 
    assign out[526] = layer_0[685] ^ layer_0[1172]; 
    assign out[527] = ~(layer_0[705] & layer_0[732]); 
    assign out[528] = layer_0[1106] ^ layer_0[215]; 
    assign out[529] = ~layer_0[1377]; 
    assign out[530] = ~(layer_0[523] ^ layer_0[415]); 
    assign out[531] = ~layer_0[1402]; 
    assign out[532] = ~(layer_0[939] ^ layer_0[1347]); 
    assign out[533] = ~(layer_0[143] ^ layer_0[1012]); 
    assign out[534] = layer_0[1216] ^ layer_0[908]; 
    assign out[535] = ~layer_0[809]; 
    assign out[536] = ~(layer_0[1483] | layer_0[718]); 
    assign out[537] = layer_0[363] | layer_0[502]; 
    assign out[538] = layer_0[892] & ~layer_0[635]; 
    assign out[539] = layer_0[216]; 
    assign out[540] = layer_0[1290]; 
    assign out[541] = layer_0[1196] & ~layer_0[1170]; 
    assign out[542] = layer_0[1466] & layer_0[476]; 
    assign out[543] = layer_0[1408] & ~layer_0[802]; 
    assign out[544] = ~layer_0[957]; 
    assign out[545] = layer_0[123] & ~layer_0[271]; 
    assign out[546] = ~layer_0[890]; 
    assign out[547] = ~(layer_0[1437] & layer_0[1413]); 
    assign out[548] = layer_0[790]; 
    assign out[549] = ~(layer_0[554] ^ layer_0[200]); 
    assign out[550] = layer_0[125]; 
    assign out[551] = layer_0[1341] & ~layer_0[1440]; 
    assign out[552] = layer_0[1098] ^ layer_0[753]; 
    assign out[553] = ~layer_0[749] | (layer_0[1162] & layer_0[749]); 
    assign out[554] = layer_0[1199] ^ layer_0[923]; 
    assign out[555] = layer_0[1291] ^ layer_0[657]; 
    assign out[556] = layer_0[1344] ^ layer_0[153]; 
    assign out[557] = ~(layer_0[1505] ^ layer_0[272]); 
    assign out[558] = ~layer_0[1163]; 
    assign out[559] = ~(layer_0[221] ^ layer_0[1382]); 
    assign out[560] = ~layer_0[768] | (layer_0[768] & layer_0[1178]); 
    assign out[561] = ~layer_0[136] | (layer_0[136] & layer_0[1260]); 
    assign out[562] = ~layer_0[937] | (layer_0[937] & layer_0[158]); 
    assign out[563] = ~(layer_0[72] ^ layer_0[659]); 
    assign out[564] = ~(layer_0[312] ^ layer_0[787]); 
    assign out[565] = layer_0[1360]; 
    assign out[566] = layer_0[1410] & layer_0[1252]; 
    assign out[567] = ~layer_0[122] | (layer_0[633] & layer_0[122]); 
    assign out[568] = layer_0[434] & layer_0[1098]; 
    assign out[569] = ~layer_0[13]; 
    assign out[570] = ~layer_0[1164]; 
    assign out[571] = ~(layer_0[1] & layer_0[703]); 
    assign out[572] = layer_0[839] ^ layer_0[1510]; 
    assign out[573] = ~layer_0[148]; 
    assign out[574] = layer_0[71]; 
    assign out[575] = ~layer_0[1479]; 
    assign out[576] = ~(layer_0[1364] ^ layer_0[981]); 
    assign out[577] = layer_0[1470] & ~layer_0[1242]; 
    assign out[578] = ~layer_0[974] | (layer_0[974] & layer_0[497]); 
    assign out[579] = ~layer_0[530]; 
    assign out[580] = layer_0[316]; 
    assign out[581] = layer_0[874] & ~layer_0[1438]; 
    assign out[582] = layer_0[495] ^ layer_0[112]; 
    assign out[583] = ~(layer_0[241] ^ layer_0[1415]); 
    assign out[584] = layer_0[1270]; 
    assign out[585] = ~(layer_0[695] ^ layer_0[1516]); 
    assign out[586] = layer_0[86]; 
    assign out[587] = ~(layer_0[737] | layer_0[1524]); 
    assign out[588] = layer_0[1361]; 
    assign out[589] = ~layer_0[1276] | (layer_0[1276] & layer_0[584]); 
    assign out[590] = layer_0[959] & layer_0[506]; 
    assign out[591] = layer_0[1207] ^ layer_0[197]; 
    assign out[592] = ~(layer_0[357] | layer_0[1373]); 
    assign out[593] = layer_0[322] & ~layer_0[1026]; 
    assign out[594] = layer_0[516] & layer_0[885]; 
    assign out[595] = layer_0[115] & ~layer_0[1129]; 
    assign out[596] = ~(layer_0[867] ^ layer_0[562]); 
    assign out[597] = layer_0[1390]; 
    assign out[598] = layer_0[654] ^ layer_0[1152]; 
    assign out[599] = ~layer_0[1379]; 
    assign out[600] = ~(layer_0[161] ^ layer_0[659]); 
    assign out[601] = layer_0[142] & ~layer_0[750]; 
    assign out[602] = layer_0[694] & layer_0[1207]; 
    assign out[603] = ~(layer_0[76] | layer_0[1307]); 
    assign out[604] = ~(layer_0[1503] | layer_0[231]); 
    assign out[605] = layer_0[879]; 
    assign out[606] = layer_0[1556] ^ layer_0[55]; 
    assign out[607] = ~layer_0[397]; 
    assign out[608] = layer_0[214] | layer_0[549]; 
    assign out[609] = layer_0[334] ^ layer_0[298]; 
    assign out[610] = layer_0[310] ^ layer_0[162]; 
    assign out[611] = ~layer_0[933]; 
    assign out[612] = ~(layer_0[598] & layer_0[900]); 
    assign out[613] = layer_0[186]; 
    assign out[614] = ~layer_0[38]; 
    assign out[615] = ~layer_0[4] | (layer_0[4] & layer_0[146]); 
    assign out[616] = layer_0[966]; 
    assign out[617] = layer_0[1266] & ~layer_0[515]; 
    assign out[618] = ~(layer_0[756] ^ layer_0[909]); 
    assign out[619] = layer_0[295] & ~layer_0[1147]; 
    assign out[620] = layer_0[1439]; 
    assign out[621] = ~layer_0[521]; 
    assign out[622] = ~(layer_0[538] ^ layer_0[717]); 
    assign out[623] = ~(layer_0[996] ^ layer_0[1113]); 
    assign out[624] = ~(layer_0[174] | layer_0[1420]); 
    assign out[625] = layer_0[536]; 
    assign out[626] = layer_0[934]; 
    assign out[627] = ~layer_0[1544]; 
    assign out[628] = layer_0[1096] ^ layer_0[784]; 
    assign out[629] = ~(layer_0[1473] ^ layer_0[207]); 
    assign out[630] = ~(layer_0[1121] ^ layer_0[607]); 
    assign out[631] = layer_0[189] & ~layer_0[1072]; 
    assign out[632] = layer_0[557]; 
    assign out[633] = ~(layer_0[1333] ^ layer_0[1535]); 
    assign out[634] = ~layer_0[1348] | (layer_0[1348] & layer_0[637]); 
    assign out[635] = layer_0[816] | layer_0[1001]; 
    assign out[636] = ~layer_0[195] | (layer_0[195] & layer_0[650]); 
    assign out[637] = ~layer_0[705]; 
    assign out[638] = ~layer_0[1472]; 
    assign out[639] = layer_0[22] ^ layer_0[1254]; 
    assign out[640] = layer_0[742] & ~layer_0[458]; 
    assign out[641] = layer_0[97]; 
    assign out[642] = layer_0[506] ^ layer_0[1179]; 
    assign out[643] = layer_0[1249] ^ layer_0[376]; 
    assign out[644] = layer_0[414] & layer_0[863]; 
    assign out[645] = layer_0[640] ^ layer_0[1067]; 
    assign out[646] = layer_0[638]; 
    assign out[647] = ~(layer_0[26] ^ layer_0[144]); 
    assign out[648] = ~layer_0[251]; 
    assign out[649] = ~(layer_0[399] ^ layer_0[83]); 
    assign out[650] = layer_0[811] & ~layer_0[1126]; 
    assign out[651] = ~layer_0[1506] | (layer_0[1506] & layer_0[1295]); 
    assign out[652] = layer_0[408] ^ layer_0[1232]; 
    assign out[653] = ~(layer_0[0] ^ layer_0[1228]); 
    assign out[654] = ~layer_0[867] | (layer_0[789] & layer_0[867]); 
    assign out[655] = layer_0[640] | layer_0[1122]; 
    assign out[656] = ~(layer_0[60] & layer_0[784]); 
    assign out[657] = ~(layer_0[56] ^ layer_0[230]); 
    assign out[658] = ~(layer_0[922] | layer_0[303]); 
    assign out[659] = ~(layer_0[263] ^ layer_0[1547]); 
    assign out[660] = layer_0[1109]; 
    assign out[661] = layer_0[1243]; 
    assign out[662] = layer_0[11] & ~layer_0[393]; 
    assign out[663] = layer_0[230] ^ layer_0[1036]; 
    assign out[664] = layer_0[1061] ^ layer_0[1366]; 
    assign out[665] = layer_0[1570]; 
    assign out[666] = ~layer_0[405]; 
    assign out[667] = layer_0[1247] | layer_0[634]; 
    assign out[668] = ~layer_0[1552] | (layer_0[514] & layer_0[1552]); 
    assign out[669] = layer_0[777] & layer_0[270]; 
    assign out[670] = layer_0[1407]; 
    assign out[671] = layer_0[971] & ~layer_0[208]; 
    assign out[672] = ~layer_0[1268]; 
    assign out[673] = ~(layer_0[992] ^ layer_0[150]); 
    assign out[674] = ~(layer_0[1041] | layer_0[1162]); 
    assign out[675] = layer_0[1285] ^ layer_0[1268]; 
    assign out[676] = ~layer_0[293]; 
    assign out[677] = ~(layer_0[369] ^ layer_0[845]); 
    assign out[678] = ~(layer_0[1332] ^ layer_0[198]); 
    assign out[679] = layer_0[1090] ^ layer_0[80]; 
    assign out[680] = layer_0[913] & ~layer_0[827]; 
    assign out[681] = layer_0[1062] ^ layer_0[165]; 
    assign out[682] = ~(layer_0[1518] | layer_0[1410]); 
    assign out[683] = ~layer_0[949]; 
    assign out[684] = layer_0[317] ^ layer_0[1202]; 
    assign out[685] = ~layer_0[644]; 
    assign out[686] = ~(layer_0[706] ^ layer_0[998]); 
    assign out[687] = layer_0[509] ^ layer_0[1589]; 
    assign out[688] = layer_0[1378] ^ layer_0[1430]; 
    assign out[689] = layer_0[1242] ^ layer_0[1353]; 
    assign out[690] = ~(layer_0[1328] ^ layer_0[991]); 
    assign out[691] = ~(layer_0[60] ^ layer_0[940]); 
    assign out[692] = layer_0[779] ^ layer_0[997]; 
    assign out[693] = ~layer_0[1368] | (layer_0[758] & layer_0[1368]); 
    assign out[694] = ~(layer_0[275] ^ layer_0[1137]); 
    assign out[695] = ~layer_0[1456] | (layer_0[380] & layer_0[1456]); 
    assign out[696] = layer_0[1480] ^ layer_0[1521]; 
    assign out[697] = ~(layer_0[81] & layer_0[406]); 
    assign out[698] = layer_0[90] ^ layer_0[169]; 
    assign out[699] = ~(layer_0[247] ^ layer_0[222]); 
    assign out[700] = layer_0[176] ^ layer_0[1214]; 
    assign out[701] = ~(layer_0[1422] ^ layer_0[1512]); 
    assign out[702] = ~layer_0[249] | (layer_0[1399] & layer_0[249]); 
    assign out[703] = layer_0[770] ^ layer_0[1464]; 
    assign out[704] = ~layer_0[28] | (layer_0[286] & layer_0[28]); 
    assign out[705] = layer_0[1269] ^ layer_0[1200]; 
    assign out[706] = layer_0[1226] ^ layer_0[268]; 
    assign out[707] = ~(layer_0[63] ^ layer_0[977]); 
    assign out[708] = layer_0[566] ^ layer_0[938]; 
    assign out[709] = layer_0[1163]; 
    assign out[710] = ~layer_0[1028] | (layer_0[564] & layer_0[1028]); 
    assign out[711] = layer_0[755] | layer_0[754]; 
    assign out[712] = layer_0[1573] ^ layer_0[726]; 
    assign out[713] = layer_0[1320] ^ layer_0[1497]; 
    assign out[714] = layer_0[737]; 
    assign out[715] = layer_0[128]; 
    assign out[716] = ~(layer_0[1523] ^ layer_0[29]); 
    assign out[717] = layer_0[638] ^ layer_0[215]; 
    assign out[718] = ~layer_0[1167]; 
    assign out[719] = ~layer_0[969]; 
    assign out[720] = layer_0[748]; 
    assign out[721] = ~(layer_0[910] ^ layer_0[412]); 
    assign out[722] = ~layer_0[386]; 
    assign out[723] = layer_0[147] ^ layer_0[547]; 
    assign out[724] = ~layer_0[1279]; 
    assign out[725] = ~(layer_0[1066] & layer_0[180]); 
    assign out[726] = layer_0[709]; 
    assign out[727] = ~(layer_0[1442] ^ layer_0[1346]); 
    assign out[728] = layer_0[826]; 
    assign out[729] = layer_0[1488]; 
    assign out[730] = ~layer_0[1311] | (layer_0[1141] & layer_0[1311]); 
    assign out[731] = layer_0[335] ^ layer_0[704]; 
    assign out[732] = ~(layer_0[266] ^ layer_0[652]); 
    assign out[733] = layer_0[533] & ~layer_0[895]; 
    assign out[734] = ~layer_0[738]; 
    assign out[735] = layer_0[285]; 
    assign out[736] = ~(layer_0[405] & layer_0[914]); 
    assign out[737] = layer_0[1454] & ~layer_0[688]; 
    assign out[738] = ~layer_0[1528]; 
    assign out[739] = ~(layer_0[559] ^ layer_0[236]); 
    assign out[740] = layer_0[641]; 
    assign out[741] = ~layer_0[1482] | (layer_0[697] & layer_0[1482]); 
    assign out[742] = ~layer_0[1176]; 
    assign out[743] = layer_0[468] & ~layer_0[976]; 
    assign out[744] = ~layer_0[1471] | (layer_0[239] & layer_0[1471]); 
    assign out[745] = layer_0[553] & ~layer_0[266]; 
    assign out[746] = layer_0[1225] ^ layer_0[1318]; 
    assign out[747] = ~layer_0[999]; 
    assign out[748] = ~layer_0[738]; 
    assign out[749] = ~(layer_0[1183] ^ layer_0[52]); 
    assign out[750] = layer_0[1156] ^ layer_0[1553]; 
    assign out[751] = ~(layer_0[1447] & layer_0[618]); 
    assign out[752] = layer_0[696]; 
    assign out[753] = ~(layer_0[199] ^ layer_0[1595]); 
    assign out[754] = layer_0[822] ^ layer_0[776]; 
    assign out[755] = layer_0[504] ^ layer_0[621]; 
    assign out[756] = layer_0[538] & ~layer_0[1559]; 
    assign out[757] = ~layer_0[1501] | (layer_0[929] & layer_0[1501]); 
    assign out[758] = layer_0[848] | layer_0[257]; 
    assign out[759] = layer_0[273] & layer_0[822]; 
    assign out[760] = layer_0[438] & ~layer_0[989]; 
    assign out[761] = ~layer_0[258]; 
    assign out[762] = ~(layer_0[982] & layer_0[282]); 
    assign out[763] = layer_0[1513]; 
    assign out[764] = layer_0[816] & layer_0[1331]; 
    assign out[765] = layer_0[936]; 
    assign out[766] = ~layer_0[151]; 
    assign out[767] = layer_0[550] & ~layer_0[732]; 
    assign out[768] = ~(layer_0[1177] ^ layer_0[252]); 
    assign out[769] = layer_0[1013] ^ layer_0[634]; 
    assign out[770] = layer_0[1358] & ~layer_0[1015]; 
    assign out[771] = ~(layer_0[237] | layer_0[1563]); 
    assign out[772] = ~layer_0[1388]; 
    assign out[773] = layer_0[1419] ^ layer_0[351]; 
    assign out[774] = layer_0[1173] & ~layer_0[1168]; 
    assign out[775] = ~(layer_0[1136] ^ layer_0[652]); 
    assign out[776] = ~layer_0[342]; 
    assign out[777] = ~layer_0[113]; 
    assign out[778] = ~(layer_0[805] ^ layer_0[704]); 
    assign out[779] = ~(layer_0[48] ^ layer_0[1221]); 
    assign out[780] = ~(layer_0[690] ^ layer_0[1056]); 
    assign out[781] = ~(layer_0[350] ^ layer_0[138]); 
    assign out[782] = layer_0[1107] ^ layer_0[81]; 
    assign out[783] = ~(layer_0[1590] | layer_0[496]); 
    assign out[784] = ~(layer_0[462] ^ layer_0[1301]); 
    assign out[785] = layer_0[370]; 
    assign out[786] = layer_0[472] & ~layer_0[1538]; 
    assign out[787] = layer_0[1097] & ~layer_0[1384]; 
    assign out[788] = ~(layer_0[55] ^ layer_0[89]); 
    assign out[789] = ~(layer_0[547] ^ layer_0[149]); 
    assign out[790] = layer_0[843] & ~layer_0[331]; 
    assign out[791] = layer_0[210] & ~layer_0[1283]; 
    assign out[792] = layer_0[769] & layer_0[1527]; 
    assign out[793] = layer_0[946]; 
    assign out[794] = layer_0[1353]; 
    assign out[795] = ~layer_0[863] | (layer_0[863] & layer_0[292]); 
    assign out[796] = ~(layer_0[596] | layer_0[676]); 
    assign out[797] = layer_0[725] & layer_0[152]; 
    assign out[798] = layer_0[451] ^ layer_0[1342]; 
    assign out[799] = ~(layer_0[563] | layer_0[433]); 
    assign out[800] = layer_0[775] ^ layer_0[1192]; 
    assign out[801] = ~(layer_0[699] | layer_0[347]); 
    assign out[802] = layer_0[489] & ~layer_0[478]; 
    assign out[803] = ~(layer_0[664] ^ layer_0[283]); 
    assign out[804] = layer_0[403]; 
    assign out[805] = layer_0[837] & ~layer_0[345]; 
    assign out[806] = ~layer_0[872]; 
    assign out[807] = layer_0[955]; 
    assign out[808] = layer_0[840] & ~layer_0[1076]; 
    assign out[809] = ~layer_0[1355] | (layer_0[645] & layer_0[1355]); 
    assign out[810] = ~layer_0[1484]; 
    assign out[811] = ~(layer_0[760] ^ layer_0[710]); 
    assign out[812] = layer_0[1373] & ~layer_0[519]; 
    assign out[813] = ~layer_0[624] | (layer_0[624] & layer_0[518]); 
    assign out[814] = ~(layer_0[493] ^ layer_0[1324]); 
    assign out[815] = ~layer_0[356]; 
    assign out[816] = layer_0[70]; 
    assign out[817] = layer_0[781] & layer_0[448]; 
    assign out[818] = ~(layer_0[1086] ^ layer_0[852]); 
    assign out[819] = ~(layer_0[1335] | layer_0[989]); 
    assign out[820] = layer_0[241] & ~layer_0[1193]; 
    assign out[821] = layer_0[63] ^ layer_0[1315]; 
    assign out[822] = ~(layer_0[1582] | layer_0[928]); 
    assign out[823] = layer_0[441] ^ layer_0[312]; 
    assign out[824] = layer_0[316]; 
    assign out[825] = layer_0[866] & ~layer_0[299]; 
    assign out[826] = ~layer_0[849] | (layer_0[849] & layer_0[954]); 
    assign out[827] = layer_0[1504]; 
    assign out[828] = layer_0[1133] & ~layer_0[570]; 
    assign out[829] = layer_0[297] ^ layer_0[344]; 
    assign out[830] = layer_0[163] & ~layer_0[1161]; 
    assign out[831] = layer_0[5] ^ layer_0[543]; 
    assign out[832] = ~(layer_0[313] | layer_0[53]); 
    assign out[833] = ~(layer_0[87] & layer_0[762]); 
    assign out[834] = layer_0[1544] & layer_0[290]; 
    assign out[835] = ~(layer_0[1567] | layer_0[870]); 
    assign out[836] = layer_0[780] & layer_0[990]; 
    assign out[837] = ~layer_0[349]; 
    assign out[838] = layer_0[799] & layer_0[604]; 
    assign out[839] = ~layer_0[218] | (layer_0[218] & layer_0[528]); 
    assign out[840] = layer_0[1131]; 
    assign out[841] = layer_0[12] | layer_0[1576]; 
    assign out[842] = layer_0[336] ^ layer_0[1406]; 
    assign out[843] = ~(layer_0[1345] ^ layer_0[1125]); 
    assign out[844] = layer_0[869] & ~layer_0[807]; 
    assign out[845] = ~layer_0[849] | (layer_0[1566] & layer_0[849]); 
    assign out[846] = layer_0[515]; 
    assign out[847] = ~layer_0[864] | (layer_0[864] & layer_0[828]); 
    assign out[848] = ~layer_0[1112] | (layer_0[1112] & layer_0[431]); 
    assign out[849] = ~(layer_0[170] | layer_0[798]); 
    assign out[850] = layer_0[951]; 
    assign out[851] = layer_0[47] ^ layer_0[1088]; 
    assign out[852] = ~(layer_0[338] ^ layer_0[1362]); 
    assign out[853] = ~(layer_0[423] ^ layer_0[333]); 
    assign out[854] = ~(layer_0[1250] | layer_0[1520]); 
    assign out[855] = layer_0[278] | layer_0[625]; 
    assign out[856] = ~layer_0[891] | (layer_0[36] & layer_0[891]); 
    assign out[857] = layer_0[511] & ~layer_0[228]; 
    assign out[858] = ~(layer_0[353] ^ layer_0[223]); 
    assign out[859] = ~(layer_0[1436] | layer_0[966]); 
    assign out[860] = layer_0[436] & ~layer_0[853]; 
    assign out[861] = layer_0[394] | layer_0[1376]; 
    assign out[862] = ~(layer_0[498] ^ layer_0[1135]); 
    assign out[863] = layer_0[1356]; 
    assign out[864] = layer_0[740] & layer_0[392]; 
    assign out[865] = layer_0[1059] & ~layer_0[907]; 
    assign out[866] = ~layer_0[642]; 
    assign out[867] = ~(layer_0[994] & layer_0[1053]); 
    assign out[868] = ~layer_0[1095] | (layer_0[132] & layer_0[1095]); 
    assign out[869] = layer_0[1598]; 
    assign out[870] = layer_0[1338] & ~layer_0[1519]; 
    assign out[871] = ~layer_0[383]; 
    assign out[872] = ~(layer_0[1183] ^ layer_0[1512]); 
    assign out[873] = layer_0[540] & ~layer_0[399]; 
    assign out[874] = ~layer_0[1071] | (layer_0[1071] & layer_0[1424]); 
    assign out[875] = layer_0[1447]; 
    assign out[876] = ~layer_0[510] | (layer_0[1081] & layer_0[510]); 
    assign out[877] = ~(layer_0[328] ^ layer_0[701]); 
    assign out[878] = layer_0[656]; 
    assign out[879] = ~layer_0[390] | (layer_0[390] & layer_0[683]); 
    assign out[880] = layer_0[922]; 
    assign out[881] = ~(layer_0[421] ^ layer_0[875]); 
    assign out[882] = ~(layer_0[1099] | layer_0[1517]); 
    assign out[883] = layer_0[190] & ~layer_0[220]; 
    assign out[884] = ~(layer_0[1590] | layer_0[128]); 
    assign out[885] = layer_0[1441] ^ layer_0[1548]; 
    assign out[886] = ~(layer_0[786] ^ layer_0[613]); 
    assign out[887] = ~layer_0[911]; 
    assign out[888] = ~(layer_0[1083] | layer_0[524]); 
    assign out[889] = ~(layer_0[1238] | layer_0[164]); 
    assign out[890] = ~layer_0[1453]; 
    assign out[891] = ~(layer_0[289] ^ layer_0[8]); 
    assign out[892] = layer_0[1186] ^ layer_0[296]; 
    assign out[893] = ~layer_0[99] | (layer_0[99] & layer_0[958]); 
    assign out[894] = layer_0[660] ^ layer_0[1149]; 
    assign out[895] = ~(layer_0[20] | layer_0[1093]); 
    assign out[896] = ~(layer_0[831] ^ layer_0[964]); 
    assign out[897] = ~(layer_0[1526] & layer_0[1386]); 
    assign out[898] = ~(layer_0[599] | layer_0[382]); 
    assign out[899] = ~(layer_0[1038] | layer_0[747]); 
    assign out[900] = layer_0[327] ^ layer_0[1263]; 
    assign out[901] = ~layer_0[1100]; 
    assign out[902] = layer_0[721]; 
    assign out[903] = layer_0[592]; 
    assign out[904] = layer_0[1199] ^ layer_0[225]; 
    assign out[905] = layer_0[730] | layer_0[1099]; 
    assign out[906] = ~layer_0[361]; 
    assign out[907] = ~(layer_0[102] | layer_0[407]); 
    assign out[908] = ~layer_0[38]; 
    assign out[909] = layer_0[1469] & ~layer_0[1376]; 
    assign out[910] = ~(layer_0[621] & layer_0[1184]); 
    assign out[911] = layer_0[127]; 
    assign out[912] = ~layer_0[32]; 
    assign out[913] = ~(layer_0[1018] ^ layer_0[1239]); 
    assign out[914] = layer_0[1465] ^ layer_0[629]; 
    assign out[915] = layer_0[1315] & ~layer_0[728]; 
    assign out[916] = ~(layer_0[1316] & layer_0[866]); 
    assign out[917] = ~(layer_0[823] ^ layer_0[1020]); 
    assign out[918] = ~layer_0[211]; 
    assign out[919] = ~(layer_0[471] ^ layer_0[631]); 
    assign out[920] = layer_0[719] ^ layer_0[172]; 
    assign out[921] = layer_0[1011] & ~layer_0[98]; 
    assign out[922] = ~(layer_0[527] ^ layer_0[1385]); 
    assign out[923] = layer_0[142]; 
    assign out[924] = layer_0[513]; 
    assign out[925] = layer_0[757] & layer_0[1198]; 
    assign out[926] = layer_0[988] & layer_0[46]; 
    assign out[927] = layer_0[116] & layer_0[699]; 
    assign out[928] = ~(layer_0[286] | layer_0[3]); 
    assign out[929] = ~(layer_0[533] ^ layer_0[1571]); 
    assign out[930] = layer_0[324]; 
    assign out[931] = layer_0[473] ^ layer_0[156]; 
    assign out[932] = layer_0[864]; 
    assign out[933] = ~(layer_0[885] ^ layer_0[673]); 
    assign out[934] = layer_0[1517]; 
    assign out[935] = layer_0[213] & ~layer_0[829]; 
    assign out[936] = ~layer_0[346] | (layer_0[346] & layer_0[258]); 
    assign out[937] = layer_0[896] ^ layer_0[858]; 
    assign out[938] = ~layer_0[1053]; 
    assign out[939] = ~(layer_0[1186] ^ layer_0[280]); 
    assign out[940] = ~(layer_0[617] | layer_0[260]); 
    assign out[941] = layer_0[26] ^ layer_0[1244]; 
    assign out[942] = ~layer_0[440] | (layer_0[851] & layer_0[440]); 
    assign out[943] = ~layer_0[1241]; 
    assign out[944] = layer_0[1281] ^ layer_0[553]; 
    assign out[945] = layer_0[1194] & ~layer_0[1565]; 
    assign out[946] = ~layer_0[656]; 
    assign out[947] = layer_0[1578]; 
    assign out[948] = layer_0[277] & ~layer_0[33]; 
    assign out[949] = ~(layer_0[466] ^ layer_0[317]); 
    assign out[950] = ~(layer_0[105] ^ layer_0[1246]); 
    assign out[951] = ~layer_0[51]; 
    assign out[952] = layer_0[203] & ~layer_0[1507]; 
    assign out[953] = ~layer_0[1387]; 
    assign out[954] = layer_0[459]; 
    assign out[955] = layer_0[397] & ~layer_0[333]; 
    assign out[956] = ~(layer_0[658] ^ layer_0[797]); 
    assign out[957] = layer_0[1157] & ~layer_0[1218]; 
    assign out[958] = ~(layer_0[442] ^ layer_0[107]); 
    assign out[959] = layer_0[798] & layer_0[262]; 
    assign out[960] = ~(layer_0[714] & layer_0[616]); 
    assign out[961] = ~layer_0[905]; 
    assign out[962] = layer_0[946] ^ layer_0[261]; 
    assign out[963] = layer_0[1403] | layer_0[899]; 
    assign out[964] = ~(layer_0[860] ^ layer_0[1562]); 
    assign out[965] = layer_0[34] & ~layer_0[273]; 
    assign out[966] = layer_0[1493] & layer_0[1043]; 
    assign out[967] = layer_0[363] ^ layer_0[1274]; 
    assign out[968] = layer_0[217] & ~layer_0[1300]; 
    assign out[969] = layer_0[1588] & ~layer_0[137]; 
    assign out[970] = ~(layer_0[970] | layer_0[1356]); 
    assign out[971] = ~(layer_0[542] & layer_0[944]); 
    assign out[972] = ~(layer_0[1391] | layer_0[1298]); 
    assign out[973] = layer_0[836] & layer_0[277]; 
    assign out[974] = layer_0[87] & layer_0[1275]; 
    assign out[975] = layer_0[1018]; 
    assign out[976] = ~(layer_0[734] & layer_0[1236]); 
    assign out[977] = layer_0[76] & ~layer_0[290]; 
    assign out[978] = layer_0[145] & layer_0[233]; 
    assign out[979] = ~(layer_0[1340] | layer_0[1213]); 
    assign out[980] = layer_0[546] & ~layer_0[361]; 
    assign out[981] = layer_0[311] & ~layer_0[1554]; 
    assign out[982] = ~(layer_0[532] ^ layer_0[304]); 
    assign out[983] = layer_0[1568] ^ layer_0[1334]; 
    assign out[984] = ~(layer_0[341] ^ layer_0[176]); 
    assign out[985] = layer_0[182] & ~layer_0[803]; 
    assign out[986] = ~(layer_0[386] ^ layer_0[1267]); 
    assign out[987] = ~(layer_0[709] ^ layer_0[1256]); 
    assign out[988] = layer_0[611]; 
    assign out[989] = ~(layer_0[1264] ^ layer_0[238]); 
    assign out[990] = layer_0[941] & ~layer_0[66]; 
    assign out[991] = layer_0[30] ^ layer_0[294]; 
    assign out[992] = layer_0[92] | layer_0[1502]; 
    assign out[993] = ~(layer_0[1374] ^ layer_0[1254]); 
    assign out[994] = ~(layer_0[716] ^ layer_0[479]); 
    assign out[995] = ~layer_0[599] | (layer_0[599] & layer_0[1132]); 
    assign out[996] = ~(layer_0[751] | layer_0[844]); 
    assign out[997] = layer_0[1231] & ~layer_0[1052]; 
    assign out[998] = layer_0[1599] ^ layer_0[782]; 
    assign out[999] = layer_0[379] ^ layer_0[845]; 
    assign out[1000] = ~(layer_0[917] ^ layer_0[1272]); 
    assign out[1001] = layer_0[1138]; 
    assign out[1002] = layer_0[1055]; 
    assign out[1003] = ~layer_0[724] | (layer_0[908] & layer_0[724]); 
    assign out[1004] = layer_0[579]; 
    assign out[1005] = layer_0[986] ^ layer_0[1051]; 
    assign out[1006] = layer_0[1460] & ~layer_0[582]; 
    assign out[1007] = ~layer_0[728]; 
    assign out[1008] = layer_0[1319] | layer_0[552]; 
    assign out[1009] = ~(layer_0[530] | layer_0[1259]); 
    assign out[1010] = ~(layer_0[776] ^ layer_0[920]); 
    assign out[1011] = ~(layer_0[256] ^ layer_0[559]); 
    assign out[1012] = ~layer_0[264]; 
    assign out[1013] = ~(layer_0[113] ^ layer_0[711]); 
    assign out[1014] = layer_0[578] ^ layer_0[343]; 
    assign out[1015] = ~layer_0[868]; 
    assign out[1016] = ~layer_0[1070]; 
    assign out[1017] = ~layer_0[870]; 
    assign out[1018] = layer_0[1222] ^ layer_0[435]; 
    assign out[1019] = ~(layer_0[1571] & layer_0[352]); 
    assign out[1020] = layer_0[254] | layer_0[1476]; 
    assign out[1021] = layer_0[282] | layer_0[36]; 
    assign out[1022] = ~(layer_0[632] ^ layer_0[1277]); 
    assign out[1023] = layer_0[106] ^ layer_0[1118]; 
    assign out[1024] = layer_0[1591] ^ layer_0[1453]; 
    assign out[1025] = ~(layer_0[121] ^ layer_0[544]); 
    assign out[1026] = ~(layer_0[50] | layer_0[409]); 
    assign out[1027] = layer_0[174]; 
    assign out[1028] = ~(layer_0[945] | layer_0[78]); 
    assign out[1029] = ~layer_0[1130] | (layer_0[691] & layer_0[1130]); 
    assign out[1030] = ~(layer_0[682] ^ layer_0[78]); 
    assign out[1031] = layer_0[630] & ~layer_0[402]; 
    assign out[1032] = ~(layer_0[1396] & layer_0[1396]); 
    assign out[1033] = layer_0[443] & ~layer_0[1450]; 
    assign out[1034] = layer_0[1010]; 
    assign out[1035] = layer_0[698] & layer_0[446]; 
    assign out[1036] = ~(layer_0[1451] ^ layer_0[135]); 
    assign out[1037] = ~(layer_0[768] ^ layer_0[1494]); 
    assign out[1038] = layer_0[287]; 
    assign out[1039] = layer_0[308] ^ layer_0[1197]; 
    assign out[1040] = layer_0[42] ^ layer_0[1300]; 
    assign out[1041] = ~(layer_0[325] & layer_0[608]); 
    assign out[1042] = ~layer_0[1358] | (layer_0[1358] & layer_0[1514]); 
    assign out[1043] = layer_0[219] ^ layer_0[481]; 
    assign out[1044] = layer_0[570] & layer_0[457]; 
    assign out[1045] = ~layer_0[454] | (layer_0[1471] & layer_0[454]); 
    assign out[1046] = ~(layer_0[897] ^ layer_0[1008]); 
    assign out[1047] = layer_0[460] ^ layer_0[681]; 
    assign out[1048] = ~layer_0[50]; 
    assign out[1049] = layer_0[1021]; 
    assign out[1050] = ~layer_0[1477]; 
    assign out[1051] = layer_0[1166]; 
    assign out[1052] = ~layer_0[965]; 
    assign out[1053] = ~layer_0[1513]; 
    assign out[1054] = layer_0[1225] ^ layer_0[549]; 
    assign out[1055] = layer_0[1079]; 
    assign out[1056] = layer_0[853] ^ layer_0[1174]; 
    assign out[1057] = layer_0[1000] & layer_0[675]; 
    assign out[1058] = ~(layer_0[1337] ^ layer_0[470]); 
    assign out[1059] = layer_0[519] & ~layer_0[1443]; 
    assign out[1060] = ~layer_0[1237] | (layer_0[1237] & layer_0[489]); 
    assign out[1061] = layer_0[883] | layer_0[1405]; 
    assign out[1062] = ~layer_0[586] | (layer_0[586] & layer_0[1010]); 
    assign out[1063] = layer_0[1004] ^ layer_0[1337]; 
    assign out[1064] = layer_0[765] & layer_0[561]; 
    assign out[1065] = ~(layer_0[384] ^ layer_0[548]); 
    assign out[1066] = ~(layer_0[668] ^ layer_0[749]); 
    assign out[1067] = layer_0[107]; 
    assign out[1068] = layer_0[1001] ^ layer_0[1253]; 
    assign out[1069] = layer_0[1255] & ~layer_0[427]; 
    assign out[1070] = ~(layer_0[421] ^ layer_0[560]); 
    assign out[1071] = ~layer_0[791] | (layer_0[791] & layer_0[1514]); 
    assign out[1072] = ~(layer_0[117] ^ layer_0[1150]); 
    assign out[1073] = ~layer_0[1077] | (layer_0[1077] & layer_0[635]); 
    assign out[1074] = ~layer_0[880]; 
    assign out[1075] = ~(layer_0[1461] ^ layer_0[1333]); 
    assign out[1076] = ~(layer_0[1210] ^ layer_0[1169]); 
    assign out[1077] = layer_0[1196]; 
    assign out[1078] = ~layer_0[1499] | (layer_0[335] & layer_0[1499]); 
    assign out[1079] = ~(layer_0[77] ^ layer_0[178]); 
    assign out[1080] = layer_0[766] & layer_0[119]; 
    assign out[1081] = layer_0[1087] ^ layer_0[476]; 
    assign out[1082] = ~(layer_0[366] ^ layer_0[670]); 
    assign out[1083] = ~layer_0[773]; 
    assign out[1084] = ~(layer_0[1312] ^ layer_0[927]); 
    assign out[1085] = layer_0[1586] & ~layer_0[1542]; 
    assign out[1086] = ~(layer_0[819] ^ layer_0[492]); 
    assign out[1087] = ~(layer_0[454] ^ layer_0[731]); 
    assign out[1088] = layer_0[169] ^ layer_0[846]; 
    assign out[1089] = layer_0[978] ^ layer_0[1533]; 
    assign out[1090] = ~(layer_0[792] ^ layer_0[894]); 
    assign out[1091] = layer_0[526] ^ layer_0[1208]; 
    assign out[1092] = ~(layer_0[1303] ^ layer_0[1445]); 
    assign out[1093] = ~(layer_0[296] ^ layer_0[1046]); 
    assign out[1094] = ~(layer_0[131] ^ layer_0[369]); 
    assign out[1095] = ~(layer_0[1181] ^ layer_0[1561]); 
    assign out[1096] = ~(layer_0[513] | layer_0[1508]); 
    assign out[1097] = layer_0[558] | layer_0[166]; 
    assign out[1098] = ~(layer_0[1295] | layer_0[124]); 
    assign out[1099] = ~(layer_0[298] ^ layer_0[827]); 
    assign out[1100] = ~(layer_0[1359] ^ layer_0[1435]); 
    assign out[1101] = ~(layer_0[1574] ^ layer_0[1448]); 
    assign out[1102] = layer_0[1086] | layer_0[1309]; 
    assign out[1103] = layer_0[766] & layer_0[44]; 
    assign out[1104] = layer_0[1395]; 
    assign out[1105] = ~(layer_0[778] ^ layer_0[201]); 
    assign out[1106] = ~layer_0[1433] | (layer_0[1433] & layer_0[494]); 
    assign out[1107] = ~layer_0[1564]; 
    assign out[1108] = layer_0[1062] ^ layer_0[1227]; 
    assign out[1109] = layer_0[995] ^ layer_0[16]; 
    assign out[1110] = ~layer_0[941] | (layer_0[723] & layer_0[941]); 
    assign out[1111] = ~layer_0[1188]; 
    assign out[1112] = layer_0[1078]; 
    assign out[1113] = ~(layer_0[1271] & layer_0[1354]); 
    assign out[1114] = layer_0[1391]; 
    assign out[1115] = layer_0[157] & ~layer_0[1009]; 
    assign out[1116] = layer_0[1308] & layer_0[1236]; 
    assign out[1117] = layer_0[700] ^ layer_0[683]; 
    assign out[1118] = layer_0[348]; 
    assign out[1119] = ~(layer_0[45] | layer_0[344]); 
    assign out[1120] = ~(layer_0[1415] ^ layer_0[1506]); 
    assign out[1121] = layer_0[1296] ^ layer_0[639]; 
    assign out[1122] = ~(layer_0[362] ^ layer_0[1080]); 
    assign out[1123] = layer_0[323] ^ layer_0[707]; 
    assign out[1124] = layer_0[1119]; 
    assign out[1125] = layer_0[904]; 
    assign out[1126] = layer_0[624]; 
    assign out[1127] = layer_0[588] & ~layer_0[1481]; 
    assign out[1128] = layer_0[587] & ~layer_0[612]; 
    assign out[1129] = ~(layer_0[130] ^ layer_0[1429]); 
    assign out[1130] = layer_0[1119] & ~layer_0[543]; 
    assign out[1131] = ~(layer_0[1261] ^ layer_0[24]); 
    assign out[1132] = layer_0[1367] & ~layer_0[1329]; 
    assign out[1133] = ~(layer_0[77] & layer_0[520]); 
    assign out[1134] = ~(layer_0[1221] ^ layer_0[1400]); 
    assign out[1135] = layer_0[1392] ^ layer_0[1367]; 
    assign out[1136] = layer_0[1371] | layer_0[0]; 
    assign out[1137] = layer_0[269] ^ layer_0[259]; 
    assign out[1138] = ~layer_0[39] | (layer_0[132] & layer_0[39]); 
    assign out[1139] = ~(layer_0[774] ^ layer_0[1390]); 
    assign out[1140] = ~(layer_0[958] ^ layer_0[962]); 
    assign out[1141] = ~(layer_0[1342] ^ layer_0[488]); 
    assign out[1142] = layer_0[1292] & layer_0[667]; 
    assign out[1143] = layer_0[1161] ^ layer_0[755]; 
    assign out[1144] = layer_0[1323] ^ layer_0[1452]; 
    assign out[1145] = layer_0[348] & ~layer_0[646]; 
    assign out[1146] = layer_0[1426] ^ layer_0[1246]; 
    assign out[1147] = ~(layer_0[1151] ^ layer_0[389]); 
    assign out[1148] = layer_0[465]; 
    assign out[1149] = ~layer_0[1487]; 
    assign out[1150] = layer_0[1211] & ~layer_0[1089]; 
    assign out[1151] = layer_0[1169] & ~layer_0[796]; 
    assign out[1152] = ~(layer_0[546] ^ layer_0[1224]); 
    assign out[1153] = layer_0[391] & ~layer_0[537]; 
    assign out[1154] = ~(layer_0[1032] ^ layer_0[232]); 
    assign out[1155] = ~layer_0[977]; 
    assign out[1156] = layer_0[167]; 
    assign out[1157] = layer_0[447] ^ layer_0[925]; 
    assign out[1158] = layer_0[1179]; 
    assign out[1159] = layer_0[619] ^ layer_0[1428]; 
    assign out[1160] = ~(layer_0[1042] ^ layer_0[155]); 
    assign out[1161] = ~(layer_0[903] ^ layer_0[1294]); 
    assign out[1162] = layer_0[186] & layer_0[861]; 
    assign out[1163] = ~(layer_0[304] ^ layer_0[1174]); 
    assign out[1164] = ~layer_0[1165]; 
    assign out[1165] = layer_0[293] ^ layer_0[772]; 
    assign out[1166] = layer_0[722] ^ layer_0[881]; 
    assign out[1167] = ~(layer_0[961] | layer_0[687]); 
    assign out[1168] = ~(layer_0[229] | layer_0[1148]); 
    assign out[1169] = ~(layer_0[850] ^ layer_0[1299]); 
    assign out[1170] = ~(layer_0[514] | layer_0[1123]); 
    assign out[1171] = layer_0[1143]; 
    assign out[1172] = layer_0[824] ^ layer_0[701]; 
    assign out[1173] = layer_0[285] & ~layer_0[529]; 
    assign out[1174] = ~(layer_0[1483] ^ layer_0[1190]); 
    assign out[1175] = layer_0[1055] & ~layer_0[835]; 
    assign out[1176] = ~(layer_0[330] ^ layer_0[1251]); 
    assign out[1177] = ~(layer_0[1522] | layer_0[1429]); 
    assign out[1178] = ~(layer_0[329] | layer_0[1043]); 
    assign out[1179] = ~(layer_0[202] ^ layer_0[418]); 
    assign out[1180] = layer_0[626] ^ layer_0[284]; 
    assign out[1181] = layer_0[931] ^ layer_0[1075]; 
    assign out[1182] = layer_0[387] ^ layer_0[800]; 
    assign out[1183] = ~layer_0[1397] | (layer_0[1397] & layer_0[1523]); 
    assign out[1184] = ~layer_0[375] | (layer_0[375] & layer_0[497]); 
    assign out[1185] = ~(layer_0[1296] ^ layer_0[575]); 
    assign out[1186] = layer_0[214] ^ layer_0[1496]; 
    assign out[1187] = ~layer_0[586]; 
    assign out[1188] = layer_0[1316] | layer_0[856]; 
    assign out[1189] = ~(layer_0[1058] & layer_0[818]); 
    assign out[1190] = layer_0[1194]; 
    assign out[1191] = ~layer_0[675] | (layer_0[675] & layer_0[193]); 
    assign out[1192] = ~(layer_0[1546] ^ layer_0[752]); 
    assign out[1193] = ~(layer_0[59] | layer_0[577]); 
    assign out[1194] = layer_0[536] & ~layer_0[1343]; 
    assign out[1195] = ~layer_0[1293]; 
    assign out[1196] = ~(layer_0[181] | layer_0[1313]); 
    assign out[1197] = ~(layer_0[540] ^ layer_0[1212]); 
    assign out[1198] = ~layer_0[1498] | (layer_0[1498] & layer_0[591]); 
    assign out[1199] = layer_0[1386] & ~layer_0[1566]; 
    assign out[1200] = ~(layer_0[939] | layer_0[59]); 
    assign out[1201] = ~(layer_0[263] | layer_0[684]); 
    assign out[1202] = ~layer_0[692]; 
    assign out[1203] = ~layer_0[743]; 
    assign out[1204] = layer_0[111] ^ layer_0[177]; 
    assign out[1205] = ~(layer_0[567] ^ layer_0[770]); 
    assign out[1206] = ~(layer_0[140] ^ layer_0[346]); 
    assign out[1207] = ~(layer_0[815] ^ layer_0[1455]); 
    assign out[1208] = layer_0[173] | layer_0[907]; 
    assign out[1209] = layer_0[914] & ~layer_0[1598]; 
    assign out[1210] = layer_0[1579] & layer_0[28]; 
    assign out[1211] = layer_0[920] & layer_0[257]; 
    assign out[1212] = ~(layer_0[306] ^ layer_0[935]); 
    assign out[1213] = layer_0[1103] & ~layer_0[756]; 
    assign out[1214] = ~layer_0[686] | (layer_0[736] & layer_0[686]); 
    assign out[1215] = ~(layer_0[842] | layer_0[499]); 
    assign out[1216] = ~(layer_0[1350] & layer_0[1301]); 
    assign out[1217] = ~(layer_0[663] | layer_0[1400]); 
    assign out[1218] = layer_0[1297] & ~layer_0[102]; 
    assign out[1219] = layer_0[1394] & layer_0[1151]; 
    assign out[1220] = ~(layer_0[288] ^ layer_0[1084]); 
    assign out[1221] = ~(layer_0[1477] | layer_0[544]); 
    assign out[1222] = ~(layer_0[636] ^ layer_0[237]); 
    assign out[1223] = ~(layer_0[1149] & layer_0[1592]); 
    assign out[1224] = layer_0[1231] ^ layer_0[356]; 
    assign out[1225] = ~(layer_0[1002] ^ layer_0[463]); 
    assign out[1226] = layer_0[490] & layer_0[1482]; 
    assign out[1227] = ~(layer_0[1108] ^ layer_0[91]); 
    assign out[1228] = layer_0[82]; 
    assign out[1229] = ~layer_0[1229] | (layer_0[1085] & layer_0[1229]); 
    assign out[1230] = ~(layer_0[842] | layer_0[956]); 
    assign out[1231] = layer_0[825]; 
    assign out[1232] = ~layer_0[392]; 
    assign out[1233] = ~(layer_0[679] ^ layer_0[491]); 
    assign out[1234] = ~(layer_0[1064] | layer_0[682]); 
    assign out[1235] = layer_0[881] ^ layer_0[1251]; 
    assign out[1236] = layer_0[851] ^ layer_0[931]; 
    assign out[1237] = layer_0[193]; 
    assign out[1238] = ~(layer_0[1393] & layer_0[1542]); 
    assign out[1239] = layer_0[1013] & ~layer_0[279]; 
    assign out[1240] = layer_0[1110] | layer_0[1233]; 
    assign out[1241] = layer_0[522]; 
    assign out[1242] = ~layer_0[535] | (layer_0[535] & layer_0[467]); 
    assign out[1243] = layer_0[1021] & ~layer_0[152]; 
    assign out[1244] = layer_0[1244] ^ layer_0[329]; 
    assign out[1245] = layer_0[935] & ~layer_0[615]; 
    assign out[1246] = layer_0[74] & layer_0[1115]; 
    assign out[1247] = layer_0[62] ^ layer_0[824]; 
    assign out[1248] = layer_0[661] & layer_0[919]; 
    assign out[1249] = layer_0[1475] & layer_0[1304]; 
    assign out[1250] = layer_0[1576]; 
    assign out[1251] = layer_0[159] & ~layer_0[1278]; 
    assign out[1252] = layer_0[1427] & ~layer_0[1224]; 
    assign out[1253] = ~(layer_0[1222] ^ layer_0[187]); 
    assign out[1254] = ~(layer_0[1154] & layer_0[1201]); 
    assign out[1255] = ~(layer_0[1282] ^ layer_0[1458]); 
    assign out[1256] = layer_0[1444] & layer_0[480]; 
    assign out[1257] = ~layer_0[1375]; 
    assign out[1258] = ~(layer_0[1310] | layer_0[921]); 
    assign out[1259] = layer_0[72] ^ layer_0[199]; 
    assign out[1260] = ~layer_0[576] | (layer_0[576] & layer_0[930]); 
    assign out[1261] = ~layer_0[1031] | (layer_0[191] & layer_0[1031]); 
    assign out[1262] = ~(layer_0[68] ^ layer_0[485]); 
    assign out[1263] = ~(layer_0[1101] ^ layer_0[274]); 
    assign out[1264] = ~(layer_0[1409] ^ layer_0[512]); 
    assign out[1265] = ~(layer_0[471] ^ layer_0[1346]); 
    assign out[1266] = ~(layer_0[91] & layer_0[1064]); 
    assign out[1267] = ~layer_0[925]; 
    assign out[1268] = ~(layer_0[720] ^ layer_0[840]); 
    assign out[1269] = layer_0[347]; 
    assign out[1270] = 1'b0; 
    assign out[1271] = 1'b0; 
    assign out[1272] = 1'b0; 
    assign out[1273] = 1'b0; 
    assign out[1274] = 1'b0; 
    assign out[1275] = 1'b0; 
    assign out[1276] = 1'b0; 
    assign out[1277] = 1'b0; 
    assign out[1278] = 1'b0; 
    assign out[1279] = 1'b0; 
    assign out[1280] = 1'b0; 
    assign out[1281] = 1'b0; 
    assign out[1282] = 1'b0; 
    assign out[1283] = 1'b0; 
    assign out[1284] = 1'b0; 
    assign out[1285] = 1'b0; 
    assign out[1286] = 1'b0; 
    assign out[1287] = 1'b0; 
    assign out[1288] = 1'b0; 
    assign out[1289] = 1'b0; 
    assign out[1290] = 1'b0; 
    assign out[1291] = 1'b0; 
    assign out[1292] = 1'b0; 
    assign out[1293] = 1'b0; 
    assign out[1294] = 1'b0; 
    assign out[1295] = 1'b0; 
    assign out[1296] = 1'b0; 
    assign out[1297] = 1'b0; 
    assign out[1298] = 1'b0; 
    assign out[1299] = 1'b0; 
    assign out[1300] = 1'b0; 
    assign out[1301] = 1'b0; 
    assign out[1302] = 1'b0; 
    assign out[1303] = 1'b0; 
    assign out[1304] = 1'b0; 
    assign out[1305] = 1'b0; 
    assign out[1306] = 1'b0; 
    assign out[1307] = 1'b0; 
    assign out[1308] = 1'b0; 
    assign out[1309] = 1'b0; 
    assign out[1310] = 1'b0; 
    assign out[1311] = 1'b0; 
    assign out[1312] = 1'b0; 
    assign out[1313] = 1'b0; 
    assign out[1314] = 1'b0; 
    assign out[1315] = 1'b0; 
    assign out[1316] = 1'b0; 
    assign out[1317] = 1'b0; 
    assign out[1318] = 1'b0; 
    assign out[1319] = 1'b0; 
    assign out[1320] = 1'b0; 
    assign out[1321] = 1'b0; 
    assign out[1322] = 1'b0; 
    assign out[1323] = 1'b0; 
    assign out[1324] = 1'b0; 
    assign out[1325] = 1'b0; 
    assign out[1326] = 1'b0; 
    assign out[1327] = 1'b0; 
    assign out[1328] = 1'b0; 
    assign out[1329] = 1'b0; 
    assign out[1330] = 1'b0; 
    assign out[1331] = 1'b0; 
    assign out[1332] = 1'b0; 
    assign out[1333] = 1'b0; 
    assign out[1334] = 1'b0; 
    assign out[1335] = 1'b0; 
    assign out[1336] = 1'b0; 
    assign out[1337] = 1'b0; 
    assign out[1338] = 1'b0; 
    assign out[1339] = 1'b0; 
    assign out[1340] = 1'b0; 
    assign out[1341] = 1'b0; 
    assign out[1342] = 1'b0; 
    assign out[1343] = 1'b0; 
    assign out[1344] = 1'b0; 
    assign out[1345] = 1'b0; 
    assign out[1346] = 1'b0; 
    assign out[1347] = 1'b0; 
    assign out[1348] = 1'b0; 
    assign out[1349] = 1'b0; 
    assign out[1350] = 1'b0; 
    assign out[1351] = 1'b0; 
    assign out[1352] = 1'b0; 
    assign out[1353] = 1'b0; 
    assign out[1354] = 1'b0; 
    assign out[1355] = 1'b0; 
    assign out[1356] = 1'b0; 
    assign out[1357] = 1'b0; 
    assign out[1358] = 1'b0; 
    assign out[1359] = 1'b0; 
    assign out[1360] = 1'b0; 
    assign out[1361] = 1'b0; 
    assign out[1362] = 1'b0; 
    assign out[1363] = 1'b0; 
    assign out[1364] = 1'b0; 
    assign out[1365] = 1'b0; 
    assign out[1366] = 1'b0; 
    assign out[1367] = 1'b0; 
    assign out[1368] = 1'b0; 
    assign out[1369] = 1'b0; 
    assign out[1370] = 1'b0; 
    assign out[1371] = 1'b0; 
    assign out[1372] = 1'b0; 
    assign out[1373] = 1'b0; 
    assign out[1374] = 1'b0; 
    assign out[1375] = 1'b0; 
    assign out[1376] = 1'b0; 
    assign out[1377] = 1'b0; 
    assign out[1378] = 1'b0; 
    assign out[1379] = 1'b0; 
    assign out[1380] = 1'b0; 
    assign out[1381] = 1'b0; 
    assign out[1382] = 1'b0; 
    assign out[1383] = 1'b0; 
    assign out[1384] = 1'b0; 
    assign out[1385] = 1'b0; 
    assign out[1386] = 1'b0; 
    assign out[1387] = 1'b0; 
    assign out[1388] = 1'b0; 
    assign out[1389] = 1'b0; 
    assign out[1390] = 1'b0; 
    assign out[1391] = 1'b0; 
    assign out[1392] = 1'b0; 
    assign out[1393] = 1'b0; 
    assign out[1394] = 1'b0; 
    assign out[1395] = 1'b0; 
    assign out[1396] = 1'b0; 
    assign out[1397] = 1'b0; 
    assign out[1398] = 1'b0; 
    assign out[1399] = 1'b0; 
    assign out[1400] = 1'b0; 
    assign out[1401] = 1'b0; 
    assign out[1402] = 1'b0; 
    assign out[1403] = 1'b0; 
    assign out[1404] = 1'b0; 
    assign out[1405] = 1'b0; 
    assign out[1406] = 1'b0; 
    assign out[1407] = 1'b0; 
    assign out[1408] = 1'b0; 
    assign out[1409] = 1'b0; 
    assign out[1410] = 1'b0; 
    assign out[1411] = 1'b0; 
    assign out[1412] = 1'b0; 
    assign out[1413] = 1'b0; 
    assign out[1414] = 1'b0; 
    assign out[1415] = 1'b0; 
    assign out[1416] = 1'b0; 
    assign out[1417] = 1'b0; 
    assign out[1418] = 1'b0; 
    assign out[1419] = 1'b0; 
    assign out[1420] = 1'b0; 
    assign out[1421] = 1'b0; 
    assign out[1422] = 1'b0; 
    assign out[1423] = 1'b0; 
    assign out[1424] = 1'b0; 
    assign out[1425] = 1'b0; 
    assign out[1426] = 1'b0; 
    assign out[1427] = 1'b0; 
    assign out[1428] = 1'b0; 
    assign out[1429] = 1'b0; 
    assign out[1430] = 1'b0; 
    assign out[1431] = 1'b0; 
    assign out[1432] = 1'b0; 
    assign out[1433] = 1'b0; 
    assign out[1434] = 1'b0; 
    assign out[1435] = 1'b0; 
    assign out[1436] = 1'b0; 
    assign out[1437] = 1'b0; 
    assign out[1438] = 1'b0; 
    assign out[1439] = 1'b0; 
    assign out[1440] = 1'b0; 
    assign out[1441] = 1'b0; 
    assign out[1442] = 1'b0; 
    assign out[1443] = 1'b0; 
    assign out[1444] = 1'b0; 
    assign out[1445] = 1'b0; 
    assign out[1446] = 1'b0; 
    assign out[1447] = 1'b0; 
    assign out[1448] = 1'b0; 
    assign out[1449] = 1'b0; 
    assign out[1450] = 1'b0; 
    assign out[1451] = 1'b0; 
    assign out[1452] = 1'b0; 
    assign out[1453] = 1'b0; 
    assign out[1454] = 1'b0; 
    assign out[1455] = 1'b0; 
    assign out[1456] = 1'b0; 
    assign out[1457] = 1'b0; 
    assign out[1458] = 1'b0; 
    assign out[1459] = 1'b0; 
    assign out[1460] = 1'b0; 
    assign out[1461] = 1'b0; 
    assign out[1462] = 1'b0; 
    assign out[1463] = 1'b0; 
    assign out[1464] = 1'b0; 
    assign out[1465] = 1'b0; 
    assign out[1466] = 1'b0; 
    assign out[1467] = 1'b0; 
    assign out[1468] = 1'b0; 
    assign out[1469] = 1'b0; 
    assign out[1470] = 1'b0; 
    assign out[1471] = 1'b0; 
    assign out[1472] = 1'b0; 
    assign out[1473] = 1'b0; 
    assign out[1474] = 1'b0; 
    assign out[1475] = 1'b0; 
    assign out[1476] = 1'b0; 
    assign out[1477] = 1'b0; 
    assign out[1478] = 1'b0; 
    assign out[1479] = 1'b0; 
    assign out[1480] = 1'b0; 
    assign out[1481] = 1'b0; 
    assign out[1482] = 1'b0; 
    assign out[1483] = 1'b0; 
    assign out[1484] = 1'b0; 
    assign out[1485] = 1'b0; 
    assign out[1486] = 1'b0; 
    assign out[1487] = 1'b0; 
    assign out[1488] = 1'b0; 
    assign out[1489] = 1'b0; 
    assign out[1490] = 1'b0; 
    assign out[1491] = 1'b0; 
    assign out[1492] = 1'b0; 
    assign out[1493] = 1'b0; 
    assign out[1494] = 1'b0; 
    assign out[1495] = 1'b0; 
    assign out[1496] = 1'b0; 
    assign out[1497] = 1'b0; 
    assign out[1498] = 1'b0; 
    assign out[1499] = 1'b0; 
    assign out[1500] = 1'b0; 
    assign out[1501] = 1'b0; 
    assign out[1502] = 1'b0; 
    assign out[1503] = 1'b0; 
    assign out[1504] = 1'b0; 
    assign out[1505] = 1'b0; 
    assign out[1506] = 1'b0; 
    assign out[1507] = 1'b0; 
    assign out[1508] = 1'b0; 
    assign out[1509] = 1'b0; 
    assign out[1510] = 1'b0; 
    assign out[1511] = 1'b0; 
    assign out[1512] = 1'b0; 
    assign out[1513] = 1'b0; 
    assign out[1514] = 1'b0; 
    assign out[1515] = 1'b0; 
    assign out[1516] = 1'b0; 
    assign out[1517] = 1'b0; 
    assign out[1518] = 1'b0; 
    assign out[1519] = 1'b0; 
    assign out[1520] = 1'b0; 
    assign out[1521] = 1'b0; 
    assign out[1522] = 1'b0; 
    assign out[1523] = 1'b0; 
    assign out[1524] = 1'b0; 
    assign out[1525] = 1'b0; 
    assign out[1526] = 1'b0; 
    assign out[1527] = 1'b0; 
    assign out[1528] = 1'b0; 
    assign out[1529] = 1'b0; 
    assign out[1530] = 1'b0; 
    assign out[1531] = 1'b0; 
    assign out[1532] = 1'b0; 
    assign out[1533] = 1'b0; 
    assign out[1534] = 1'b0; 
    assign out[1535] = 1'b0; 
    assign out[1536] = 1'b0; 
    assign out[1537] = 1'b0; 
    assign out[1538] = 1'b0; 
    assign out[1539] = 1'b0; 
    assign out[1540] = 1'b0; 
    assign out[1541] = 1'b0; 
    assign out[1542] = 1'b0; 
    assign out[1543] = 1'b0; 
    assign out[1544] = 1'b0; 
    assign out[1545] = 1'b0; 
    assign out[1546] = 1'b0; 
    assign out[1547] = 1'b0; 
    assign out[1548] = 1'b0; 
    assign out[1549] = 1'b0; 
    assign out[1550] = 1'b0; 
    assign out[1551] = 1'b0; 
    assign out[1552] = 1'b0; 
    assign out[1553] = 1'b0; 
    assign out[1554] = 1'b0; 
    assign out[1555] = 1'b0; 
    assign out[1556] = 1'b0; 
    assign out[1557] = 1'b0; 
    assign out[1558] = 1'b0; 
    assign out[1559] = 1'b0; 
    assign out[1560] = 1'b0; 
    assign out[1561] = 1'b0; 
    assign out[1562] = 1'b0; 
    assign out[1563] = 1'b0; 
    assign out[1564] = 1'b0; 
    assign out[1565] = 1'b0; 
    assign out[1566] = 1'b0; 
    assign out[1567] = 1'b0; 
    assign out[1568] = 1'b0; 
    assign out[1569] = 1'b0; 
    assign out[1570] = 1'b0; 
    assign out[1571] = 1'b0; 
    assign out[1572] = 1'b0; 
    assign out[1573] = 1'b0; 
    assign out[1574] = 1'b0; 
    assign out[1575] = 1'b0; 
    assign out[1576] = 1'b0; 
    assign out[1577] = 1'b0; 
    assign out[1578] = 1'b0; 
    assign out[1579] = 1'b0; 
    assign out[1580] = 1'b0; 
    assign out[1581] = 1'b0; 
    assign out[1582] = 1'b0; 
    assign out[1583] = 1'b0; 
    assign out[1584] = 1'b0; 
    assign out[1585] = 1'b0; 
    assign out[1586] = 1'b0; 
    assign out[1587] = 1'b0; 
    assign out[1588] = 1'b0; 
    assign out[1589] = 1'b0; 
    assign out[1590] = 1'b0; 
    assign out[1591] = 1'b0; 
    assign out[1592] = 1'b0; 
    assign out[1593] = 1'b0; 
    assign out[1594] = 1'b0; 
    assign out[1595] = 1'b0; 
    assign out[1596] = 1'b0; 
    assign out[1597] = 1'b0; 
    assign out[1598] = 1'b0; 
    assign out[1599] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[1269:0] = out[1269:0];
    // assign categories[126:0] = out[126:0];
    // assign categories[253:127] = out[286:160];
    // assign categories[380:254] = out[446:320];
    // assign categories[507:381] = out[606:480];
    // assign categories[634:508] = out[766:640];
    // assign categories[761:635] = out[926:800];
    // assign categories[888:762] = out[1086:960];
    // assign categories[1015:889] = out[1246:1120];
    // assign categories[1142:1016] = out[1406:1280];
    // assign categories[1269:1143] = out[1566:1440];

endmodule
