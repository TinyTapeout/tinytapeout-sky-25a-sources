magic
tech sky130A
magscale 1 2
timestamp 1757128580
<< nwell >>
rect -1809 -397 1809 397
<< mvpmos >>
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
<< mvpdiff >>
rect -1609 88 -1551 100
rect -1609 -88 -1597 88
rect -1563 -88 -1551 88
rect -1609 -100 -1551 -88
rect -1451 88 -1393 100
rect -1451 -88 -1439 88
rect -1405 -88 -1393 88
rect -1451 -100 -1393 -88
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
rect 1393 88 1451 100
rect 1393 -88 1405 88
rect 1439 -88 1451 88
rect 1393 -100 1451 -88
rect 1551 88 1609 100
rect 1551 -88 1563 88
rect 1597 -88 1609 88
rect 1551 -100 1609 -88
<< mvpdiffc >>
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
<< mvnsubdiff >>
rect -1743 319 1743 331
rect -1743 285 -1635 319
rect 1635 285 1743 319
rect -1743 273 1743 285
rect -1743 223 -1685 273
rect -1743 -223 -1731 223
rect -1697 -223 -1685 223
rect 1685 223 1743 273
rect -1743 -273 -1685 -223
rect 1685 -223 1697 223
rect 1731 -223 1743 223
rect 1685 -273 1743 -223
rect -1743 -285 1743 -273
rect -1743 -319 -1635 -285
rect 1635 -319 1743 -285
rect -1743 -331 1743 -319
<< mvnsubdiffcont >>
rect -1635 285 1635 319
rect -1731 -223 -1697 223
rect 1697 -223 1731 223
rect -1635 -319 1635 -285
<< poly >>
rect -1551 181 -1451 197
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1551 100 -1451 147
rect -1393 181 -1293 197
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1393 100 -1293 147
rect -1235 181 -1135 197
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1235 100 -1135 147
rect -1077 181 -977 197
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -1077 100 -977 147
rect -919 181 -819 197
rect -919 147 -903 181
rect -835 147 -819 181
rect -919 100 -819 147
rect -761 181 -661 197
rect -761 147 -745 181
rect -677 147 -661 181
rect -761 100 -661 147
rect -603 181 -503 197
rect -603 147 -587 181
rect -519 147 -503 181
rect -603 100 -503 147
rect -445 181 -345 197
rect -445 147 -429 181
rect -361 147 -345 181
rect -445 100 -345 147
rect -287 181 -187 197
rect -287 147 -271 181
rect -203 147 -187 181
rect -287 100 -187 147
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect 187 181 287 197
rect 187 147 203 181
rect 271 147 287 181
rect 187 100 287 147
rect 345 181 445 197
rect 345 147 361 181
rect 429 147 445 181
rect 345 100 445 147
rect 503 181 603 197
rect 503 147 519 181
rect 587 147 603 181
rect 503 100 603 147
rect 661 181 761 197
rect 661 147 677 181
rect 745 147 761 181
rect 661 100 761 147
rect 819 181 919 197
rect 819 147 835 181
rect 903 147 919 181
rect 819 100 919 147
rect 977 181 1077 197
rect 977 147 993 181
rect 1061 147 1077 181
rect 977 100 1077 147
rect 1135 181 1235 197
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1135 100 1235 147
rect 1293 181 1393 197
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1293 100 1393 147
rect 1451 181 1551 197
rect 1451 147 1467 181
rect 1535 147 1551 181
rect 1451 100 1551 147
rect -1551 -147 -1451 -100
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1551 -197 -1451 -181
rect -1393 -147 -1293 -100
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1393 -197 -1293 -181
rect -1235 -147 -1135 -100
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1235 -197 -1135 -181
rect -1077 -147 -977 -100
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -1077 -197 -977 -181
rect -919 -147 -819 -100
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -919 -197 -819 -181
rect -761 -147 -661 -100
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -761 -197 -661 -181
rect -603 -147 -503 -100
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -603 -197 -503 -181
rect -445 -147 -345 -100
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -445 -197 -345 -181
rect -287 -147 -187 -100
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -287 -197 -187 -181
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
rect 187 -147 287 -100
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 187 -197 287 -181
rect 345 -147 445 -100
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 345 -197 445 -181
rect 503 -147 603 -100
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 503 -197 603 -181
rect 661 -147 761 -100
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 661 -197 761 -181
rect 819 -147 919 -100
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 819 -197 919 -181
rect 977 -147 1077 -100
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 977 -197 1077 -181
rect 1135 -147 1235 -100
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1135 -197 1235 -181
rect 1293 -147 1393 -100
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1293 -197 1393 -181
rect 1451 -147 1551 -100
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect 1451 -197 1551 -181
<< polycont >>
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
<< locali >>
rect -1731 285 -1635 319
rect 1635 285 1731 319
rect -1731 223 -1697 285
rect 1697 223 1731 285
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -919 147 -903 181
rect -835 147 -819 181
rect -761 147 -745 181
rect -677 147 -661 181
rect -603 147 -587 181
rect -519 147 -503 181
rect -445 147 -429 181
rect -361 147 -345 181
rect -287 147 -271 181
rect -203 147 -187 181
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect 187 147 203 181
rect 271 147 287 181
rect 345 147 361 181
rect 429 147 445 181
rect 503 147 519 181
rect 587 147 603 181
rect 661 147 677 181
rect 745 147 761 181
rect 819 147 835 181
rect 903 147 919 181
rect 977 147 993 181
rect 1061 147 1077 181
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1451 147 1467 181
rect 1535 147 1551 181
rect -1597 88 -1563 104
rect -1597 -104 -1563 -88
rect -1439 88 -1405 104
rect -1439 -104 -1405 -88
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect 1405 88 1439 104
rect 1405 -104 1439 -88
rect 1563 88 1597 104
rect 1563 -104 1597 -88
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect -1731 -285 -1697 -223
rect 1697 -285 1731 -223
rect -1731 -319 -1635 -285
rect 1635 -319 1731 -285
<< viali >>
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
<< metal1 >>
rect -1547 181 -1455 187
rect -1547 147 -1535 181
rect -1467 147 -1455 181
rect -1547 141 -1455 147
rect -1389 181 -1297 187
rect -1389 147 -1377 181
rect -1309 147 -1297 181
rect -1389 141 -1297 147
rect -1231 181 -1139 187
rect -1231 147 -1219 181
rect -1151 147 -1139 181
rect -1231 141 -1139 147
rect -1073 181 -981 187
rect -1073 147 -1061 181
rect -993 147 -981 181
rect -1073 141 -981 147
rect -915 181 -823 187
rect -915 147 -903 181
rect -835 147 -823 181
rect -915 141 -823 147
rect -757 181 -665 187
rect -757 147 -745 181
rect -677 147 -665 181
rect -757 141 -665 147
rect -599 181 -507 187
rect -599 147 -587 181
rect -519 147 -507 181
rect -599 141 -507 147
rect -441 181 -349 187
rect -441 147 -429 181
rect -361 147 -349 181
rect -441 141 -349 147
rect -283 181 -191 187
rect -283 147 -271 181
rect -203 147 -191 181
rect -283 141 -191 147
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect 191 181 283 187
rect 191 147 203 181
rect 271 147 283 181
rect 191 141 283 147
rect 349 181 441 187
rect 349 147 361 181
rect 429 147 441 181
rect 349 141 441 147
rect 507 181 599 187
rect 507 147 519 181
rect 587 147 599 181
rect 507 141 599 147
rect 665 181 757 187
rect 665 147 677 181
rect 745 147 757 181
rect 665 141 757 147
rect 823 181 915 187
rect 823 147 835 181
rect 903 147 915 181
rect 823 141 915 147
rect 981 181 1073 187
rect 981 147 993 181
rect 1061 147 1073 181
rect 981 141 1073 147
rect 1139 181 1231 187
rect 1139 147 1151 181
rect 1219 147 1231 181
rect 1139 141 1231 147
rect 1297 181 1389 187
rect 1297 147 1309 181
rect 1377 147 1389 181
rect 1297 141 1389 147
rect 1455 181 1547 187
rect 1455 147 1467 181
rect 1535 147 1547 181
rect 1455 141 1547 147
rect -1603 88 -1557 100
rect -1603 -88 -1597 88
rect -1563 -88 -1557 88
rect -1603 -100 -1557 -88
rect -1445 88 -1399 100
rect -1445 -88 -1439 88
rect -1405 -88 -1399 88
rect -1445 -100 -1399 -88
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect 1399 88 1445 100
rect 1399 -88 1405 88
rect 1439 -88 1445 88
rect 1399 -100 1445 -88
rect 1557 88 1603 100
rect 1557 -88 1563 88
rect 1597 -88 1603 88
rect 1557 -100 1603 -88
rect -1547 -147 -1455 -141
rect -1547 -181 -1535 -147
rect -1467 -181 -1455 -147
rect -1547 -187 -1455 -181
rect -1389 -147 -1297 -141
rect -1389 -181 -1377 -147
rect -1309 -181 -1297 -147
rect -1389 -187 -1297 -181
rect -1231 -147 -1139 -141
rect -1231 -181 -1219 -147
rect -1151 -181 -1139 -147
rect -1231 -187 -1139 -181
rect -1073 -147 -981 -141
rect -1073 -181 -1061 -147
rect -993 -181 -981 -147
rect -1073 -187 -981 -181
rect -915 -147 -823 -141
rect -915 -181 -903 -147
rect -835 -181 -823 -147
rect -915 -187 -823 -181
rect -757 -147 -665 -141
rect -757 -181 -745 -147
rect -677 -181 -665 -147
rect -757 -187 -665 -181
rect -599 -147 -507 -141
rect -599 -181 -587 -147
rect -519 -181 -507 -147
rect -599 -187 -507 -181
rect -441 -147 -349 -141
rect -441 -181 -429 -147
rect -361 -181 -349 -147
rect -441 -187 -349 -181
rect -283 -147 -191 -141
rect -283 -181 -271 -147
rect -203 -181 -191 -147
rect -283 -187 -191 -181
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
rect 191 -147 283 -141
rect 191 -181 203 -147
rect 271 -181 283 -147
rect 191 -187 283 -181
rect 349 -147 441 -141
rect 349 -181 361 -147
rect 429 -181 441 -147
rect 349 -187 441 -181
rect 507 -147 599 -141
rect 507 -181 519 -147
rect 587 -181 599 -147
rect 507 -187 599 -181
rect 665 -147 757 -141
rect 665 -181 677 -147
rect 745 -181 757 -147
rect 665 -187 757 -181
rect 823 -147 915 -141
rect 823 -181 835 -147
rect 903 -181 915 -147
rect 823 -187 915 -181
rect 981 -147 1073 -141
rect 981 -181 993 -147
rect 1061 -181 1073 -147
rect 981 -187 1073 -181
rect 1139 -147 1231 -141
rect 1139 -181 1151 -147
rect 1219 -181 1231 -147
rect 1139 -187 1231 -181
rect 1297 -147 1389 -141
rect 1297 -181 1309 -147
rect 1377 -181 1389 -147
rect 1297 -187 1389 -181
rect 1455 -147 1547 -141
rect 1455 -181 1467 -147
rect 1535 -181 1547 -147
rect 1455 -187 1547 -181
<< properties >>
string FIXED_BBOX -1714 -302 1714 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
