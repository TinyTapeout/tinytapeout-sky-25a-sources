magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -1457 -1019 1457 1019
<< pmos >>
rect -1261 -800 -1061 800
rect -1003 -800 -803 800
rect -745 -800 -545 800
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
rect 545 -800 745 800
rect 803 -800 1003 800
rect 1061 -800 1261 800
<< pdiff >>
rect -1319 765 -1261 800
rect -1319 731 -1307 765
rect -1273 731 -1261 765
rect -1319 697 -1261 731
rect -1319 663 -1307 697
rect -1273 663 -1261 697
rect -1319 629 -1261 663
rect -1319 595 -1307 629
rect -1273 595 -1261 629
rect -1319 561 -1261 595
rect -1319 527 -1307 561
rect -1273 527 -1261 561
rect -1319 493 -1261 527
rect -1319 459 -1307 493
rect -1273 459 -1261 493
rect -1319 425 -1261 459
rect -1319 391 -1307 425
rect -1273 391 -1261 425
rect -1319 357 -1261 391
rect -1319 323 -1307 357
rect -1273 323 -1261 357
rect -1319 289 -1261 323
rect -1319 255 -1307 289
rect -1273 255 -1261 289
rect -1319 221 -1261 255
rect -1319 187 -1307 221
rect -1273 187 -1261 221
rect -1319 153 -1261 187
rect -1319 119 -1307 153
rect -1273 119 -1261 153
rect -1319 85 -1261 119
rect -1319 51 -1307 85
rect -1273 51 -1261 85
rect -1319 17 -1261 51
rect -1319 -17 -1307 17
rect -1273 -17 -1261 17
rect -1319 -51 -1261 -17
rect -1319 -85 -1307 -51
rect -1273 -85 -1261 -51
rect -1319 -119 -1261 -85
rect -1319 -153 -1307 -119
rect -1273 -153 -1261 -119
rect -1319 -187 -1261 -153
rect -1319 -221 -1307 -187
rect -1273 -221 -1261 -187
rect -1319 -255 -1261 -221
rect -1319 -289 -1307 -255
rect -1273 -289 -1261 -255
rect -1319 -323 -1261 -289
rect -1319 -357 -1307 -323
rect -1273 -357 -1261 -323
rect -1319 -391 -1261 -357
rect -1319 -425 -1307 -391
rect -1273 -425 -1261 -391
rect -1319 -459 -1261 -425
rect -1319 -493 -1307 -459
rect -1273 -493 -1261 -459
rect -1319 -527 -1261 -493
rect -1319 -561 -1307 -527
rect -1273 -561 -1261 -527
rect -1319 -595 -1261 -561
rect -1319 -629 -1307 -595
rect -1273 -629 -1261 -595
rect -1319 -663 -1261 -629
rect -1319 -697 -1307 -663
rect -1273 -697 -1261 -663
rect -1319 -731 -1261 -697
rect -1319 -765 -1307 -731
rect -1273 -765 -1261 -731
rect -1319 -800 -1261 -765
rect -1061 765 -1003 800
rect -1061 731 -1049 765
rect -1015 731 -1003 765
rect -1061 697 -1003 731
rect -1061 663 -1049 697
rect -1015 663 -1003 697
rect -1061 629 -1003 663
rect -1061 595 -1049 629
rect -1015 595 -1003 629
rect -1061 561 -1003 595
rect -1061 527 -1049 561
rect -1015 527 -1003 561
rect -1061 493 -1003 527
rect -1061 459 -1049 493
rect -1015 459 -1003 493
rect -1061 425 -1003 459
rect -1061 391 -1049 425
rect -1015 391 -1003 425
rect -1061 357 -1003 391
rect -1061 323 -1049 357
rect -1015 323 -1003 357
rect -1061 289 -1003 323
rect -1061 255 -1049 289
rect -1015 255 -1003 289
rect -1061 221 -1003 255
rect -1061 187 -1049 221
rect -1015 187 -1003 221
rect -1061 153 -1003 187
rect -1061 119 -1049 153
rect -1015 119 -1003 153
rect -1061 85 -1003 119
rect -1061 51 -1049 85
rect -1015 51 -1003 85
rect -1061 17 -1003 51
rect -1061 -17 -1049 17
rect -1015 -17 -1003 17
rect -1061 -51 -1003 -17
rect -1061 -85 -1049 -51
rect -1015 -85 -1003 -51
rect -1061 -119 -1003 -85
rect -1061 -153 -1049 -119
rect -1015 -153 -1003 -119
rect -1061 -187 -1003 -153
rect -1061 -221 -1049 -187
rect -1015 -221 -1003 -187
rect -1061 -255 -1003 -221
rect -1061 -289 -1049 -255
rect -1015 -289 -1003 -255
rect -1061 -323 -1003 -289
rect -1061 -357 -1049 -323
rect -1015 -357 -1003 -323
rect -1061 -391 -1003 -357
rect -1061 -425 -1049 -391
rect -1015 -425 -1003 -391
rect -1061 -459 -1003 -425
rect -1061 -493 -1049 -459
rect -1015 -493 -1003 -459
rect -1061 -527 -1003 -493
rect -1061 -561 -1049 -527
rect -1015 -561 -1003 -527
rect -1061 -595 -1003 -561
rect -1061 -629 -1049 -595
rect -1015 -629 -1003 -595
rect -1061 -663 -1003 -629
rect -1061 -697 -1049 -663
rect -1015 -697 -1003 -663
rect -1061 -731 -1003 -697
rect -1061 -765 -1049 -731
rect -1015 -765 -1003 -731
rect -1061 -800 -1003 -765
rect -803 765 -745 800
rect -803 731 -791 765
rect -757 731 -745 765
rect -803 697 -745 731
rect -803 663 -791 697
rect -757 663 -745 697
rect -803 629 -745 663
rect -803 595 -791 629
rect -757 595 -745 629
rect -803 561 -745 595
rect -803 527 -791 561
rect -757 527 -745 561
rect -803 493 -745 527
rect -803 459 -791 493
rect -757 459 -745 493
rect -803 425 -745 459
rect -803 391 -791 425
rect -757 391 -745 425
rect -803 357 -745 391
rect -803 323 -791 357
rect -757 323 -745 357
rect -803 289 -745 323
rect -803 255 -791 289
rect -757 255 -745 289
rect -803 221 -745 255
rect -803 187 -791 221
rect -757 187 -745 221
rect -803 153 -745 187
rect -803 119 -791 153
rect -757 119 -745 153
rect -803 85 -745 119
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -119 -745 -85
rect -803 -153 -791 -119
rect -757 -153 -745 -119
rect -803 -187 -745 -153
rect -803 -221 -791 -187
rect -757 -221 -745 -187
rect -803 -255 -745 -221
rect -803 -289 -791 -255
rect -757 -289 -745 -255
rect -803 -323 -745 -289
rect -803 -357 -791 -323
rect -757 -357 -745 -323
rect -803 -391 -745 -357
rect -803 -425 -791 -391
rect -757 -425 -745 -391
rect -803 -459 -745 -425
rect -803 -493 -791 -459
rect -757 -493 -745 -459
rect -803 -527 -745 -493
rect -803 -561 -791 -527
rect -757 -561 -745 -527
rect -803 -595 -745 -561
rect -803 -629 -791 -595
rect -757 -629 -745 -595
rect -803 -663 -745 -629
rect -803 -697 -791 -663
rect -757 -697 -745 -663
rect -803 -731 -745 -697
rect -803 -765 -791 -731
rect -757 -765 -745 -731
rect -803 -800 -745 -765
rect -545 765 -487 800
rect -545 731 -533 765
rect -499 731 -487 765
rect -545 697 -487 731
rect -545 663 -533 697
rect -499 663 -487 697
rect -545 629 -487 663
rect -545 595 -533 629
rect -499 595 -487 629
rect -545 561 -487 595
rect -545 527 -533 561
rect -499 527 -487 561
rect -545 493 -487 527
rect -545 459 -533 493
rect -499 459 -487 493
rect -545 425 -487 459
rect -545 391 -533 425
rect -499 391 -487 425
rect -545 357 -487 391
rect -545 323 -533 357
rect -499 323 -487 357
rect -545 289 -487 323
rect -545 255 -533 289
rect -499 255 -487 289
rect -545 221 -487 255
rect -545 187 -533 221
rect -499 187 -487 221
rect -545 153 -487 187
rect -545 119 -533 153
rect -499 119 -487 153
rect -545 85 -487 119
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -119 -487 -85
rect -545 -153 -533 -119
rect -499 -153 -487 -119
rect -545 -187 -487 -153
rect -545 -221 -533 -187
rect -499 -221 -487 -187
rect -545 -255 -487 -221
rect -545 -289 -533 -255
rect -499 -289 -487 -255
rect -545 -323 -487 -289
rect -545 -357 -533 -323
rect -499 -357 -487 -323
rect -545 -391 -487 -357
rect -545 -425 -533 -391
rect -499 -425 -487 -391
rect -545 -459 -487 -425
rect -545 -493 -533 -459
rect -499 -493 -487 -459
rect -545 -527 -487 -493
rect -545 -561 -533 -527
rect -499 -561 -487 -527
rect -545 -595 -487 -561
rect -545 -629 -533 -595
rect -499 -629 -487 -595
rect -545 -663 -487 -629
rect -545 -697 -533 -663
rect -499 -697 -487 -663
rect -545 -731 -487 -697
rect -545 -765 -533 -731
rect -499 -765 -487 -731
rect -545 -800 -487 -765
rect -287 765 -229 800
rect -287 731 -275 765
rect -241 731 -229 765
rect -287 697 -229 731
rect -287 663 -275 697
rect -241 663 -229 697
rect -287 629 -229 663
rect -287 595 -275 629
rect -241 595 -229 629
rect -287 561 -229 595
rect -287 527 -275 561
rect -241 527 -229 561
rect -287 493 -229 527
rect -287 459 -275 493
rect -241 459 -229 493
rect -287 425 -229 459
rect -287 391 -275 425
rect -241 391 -229 425
rect -287 357 -229 391
rect -287 323 -275 357
rect -241 323 -229 357
rect -287 289 -229 323
rect -287 255 -275 289
rect -241 255 -229 289
rect -287 221 -229 255
rect -287 187 -275 221
rect -241 187 -229 221
rect -287 153 -229 187
rect -287 119 -275 153
rect -241 119 -229 153
rect -287 85 -229 119
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -119 -229 -85
rect -287 -153 -275 -119
rect -241 -153 -229 -119
rect -287 -187 -229 -153
rect -287 -221 -275 -187
rect -241 -221 -229 -187
rect -287 -255 -229 -221
rect -287 -289 -275 -255
rect -241 -289 -229 -255
rect -287 -323 -229 -289
rect -287 -357 -275 -323
rect -241 -357 -229 -323
rect -287 -391 -229 -357
rect -287 -425 -275 -391
rect -241 -425 -229 -391
rect -287 -459 -229 -425
rect -287 -493 -275 -459
rect -241 -493 -229 -459
rect -287 -527 -229 -493
rect -287 -561 -275 -527
rect -241 -561 -229 -527
rect -287 -595 -229 -561
rect -287 -629 -275 -595
rect -241 -629 -229 -595
rect -287 -663 -229 -629
rect -287 -697 -275 -663
rect -241 -697 -229 -663
rect -287 -731 -229 -697
rect -287 -765 -275 -731
rect -241 -765 -229 -731
rect -287 -800 -229 -765
rect -29 765 29 800
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -800 29 -765
rect 229 765 287 800
rect 229 731 241 765
rect 275 731 287 765
rect 229 697 287 731
rect 229 663 241 697
rect 275 663 287 697
rect 229 629 287 663
rect 229 595 241 629
rect 275 595 287 629
rect 229 561 287 595
rect 229 527 241 561
rect 275 527 287 561
rect 229 493 287 527
rect 229 459 241 493
rect 275 459 287 493
rect 229 425 287 459
rect 229 391 241 425
rect 275 391 287 425
rect 229 357 287 391
rect 229 323 241 357
rect 275 323 287 357
rect 229 289 287 323
rect 229 255 241 289
rect 275 255 287 289
rect 229 221 287 255
rect 229 187 241 221
rect 275 187 287 221
rect 229 153 287 187
rect 229 119 241 153
rect 275 119 287 153
rect 229 85 287 119
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -119 287 -85
rect 229 -153 241 -119
rect 275 -153 287 -119
rect 229 -187 287 -153
rect 229 -221 241 -187
rect 275 -221 287 -187
rect 229 -255 287 -221
rect 229 -289 241 -255
rect 275 -289 287 -255
rect 229 -323 287 -289
rect 229 -357 241 -323
rect 275 -357 287 -323
rect 229 -391 287 -357
rect 229 -425 241 -391
rect 275 -425 287 -391
rect 229 -459 287 -425
rect 229 -493 241 -459
rect 275 -493 287 -459
rect 229 -527 287 -493
rect 229 -561 241 -527
rect 275 -561 287 -527
rect 229 -595 287 -561
rect 229 -629 241 -595
rect 275 -629 287 -595
rect 229 -663 287 -629
rect 229 -697 241 -663
rect 275 -697 287 -663
rect 229 -731 287 -697
rect 229 -765 241 -731
rect 275 -765 287 -731
rect 229 -800 287 -765
rect 487 765 545 800
rect 487 731 499 765
rect 533 731 545 765
rect 487 697 545 731
rect 487 663 499 697
rect 533 663 545 697
rect 487 629 545 663
rect 487 595 499 629
rect 533 595 545 629
rect 487 561 545 595
rect 487 527 499 561
rect 533 527 545 561
rect 487 493 545 527
rect 487 459 499 493
rect 533 459 545 493
rect 487 425 545 459
rect 487 391 499 425
rect 533 391 545 425
rect 487 357 545 391
rect 487 323 499 357
rect 533 323 545 357
rect 487 289 545 323
rect 487 255 499 289
rect 533 255 545 289
rect 487 221 545 255
rect 487 187 499 221
rect 533 187 545 221
rect 487 153 545 187
rect 487 119 499 153
rect 533 119 545 153
rect 487 85 545 119
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -119 545 -85
rect 487 -153 499 -119
rect 533 -153 545 -119
rect 487 -187 545 -153
rect 487 -221 499 -187
rect 533 -221 545 -187
rect 487 -255 545 -221
rect 487 -289 499 -255
rect 533 -289 545 -255
rect 487 -323 545 -289
rect 487 -357 499 -323
rect 533 -357 545 -323
rect 487 -391 545 -357
rect 487 -425 499 -391
rect 533 -425 545 -391
rect 487 -459 545 -425
rect 487 -493 499 -459
rect 533 -493 545 -459
rect 487 -527 545 -493
rect 487 -561 499 -527
rect 533 -561 545 -527
rect 487 -595 545 -561
rect 487 -629 499 -595
rect 533 -629 545 -595
rect 487 -663 545 -629
rect 487 -697 499 -663
rect 533 -697 545 -663
rect 487 -731 545 -697
rect 487 -765 499 -731
rect 533 -765 545 -731
rect 487 -800 545 -765
rect 745 765 803 800
rect 745 731 757 765
rect 791 731 803 765
rect 745 697 803 731
rect 745 663 757 697
rect 791 663 803 697
rect 745 629 803 663
rect 745 595 757 629
rect 791 595 803 629
rect 745 561 803 595
rect 745 527 757 561
rect 791 527 803 561
rect 745 493 803 527
rect 745 459 757 493
rect 791 459 803 493
rect 745 425 803 459
rect 745 391 757 425
rect 791 391 803 425
rect 745 357 803 391
rect 745 323 757 357
rect 791 323 803 357
rect 745 289 803 323
rect 745 255 757 289
rect 791 255 803 289
rect 745 221 803 255
rect 745 187 757 221
rect 791 187 803 221
rect 745 153 803 187
rect 745 119 757 153
rect 791 119 803 153
rect 745 85 803 119
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -119 803 -85
rect 745 -153 757 -119
rect 791 -153 803 -119
rect 745 -187 803 -153
rect 745 -221 757 -187
rect 791 -221 803 -187
rect 745 -255 803 -221
rect 745 -289 757 -255
rect 791 -289 803 -255
rect 745 -323 803 -289
rect 745 -357 757 -323
rect 791 -357 803 -323
rect 745 -391 803 -357
rect 745 -425 757 -391
rect 791 -425 803 -391
rect 745 -459 803 -425
rect 745 -493 757 -459
rect 791 -493 803 -459
rect 745 -527 803 -493
rect 745 -561 757 -527
rect 791 -561 803 -527
rect 745 -595 803 -561
rect 745 -629 757 -595
rect 791 -629 803 -595
rect 745 -663 803 -629
rect 745 -697 757 -663
rect 791 -697 803 -663
rect 745 -731 803 -697
rect 745 -765 757 -731
rect 791 -765 803 -731
rect 745 -800 803 -765
rect 1003 765 1061 800
rect 1003 731 1015 765
rect 1049 731 1061 765
rect 1003 697 1061 731
rect 1003 663 1015 697
rect 1049 663 1061 697
rect 1003 629 1061 663
rect 1003 595 1015 629
rect 1049 595 1061 629
rect 1003 561 1061 595
rect 1003 527 1015 561
rect 1049 527 1061 561
rect 1003 493 1061 527
rect 1003 459 1015 493
rect 1049 459 1061 493
rect 1003 425 1061 459
rect 1003 391 1015 425
rect 1049 391 1061 425
rect 1003 357 1061 391
rect 1003 323 1015 357
rect 1049 323 1061 357
rect 1003 289 1061 323
rect 1003 255 1015 289
rect 1049 255 1061 289
rect 1003 221 1061 255
rect 1003 187 1015 221
rect 1049 187 1061 221
rect 1003 153 1061 187
rect 1003 119 1015 153
rect 1049 119 1061 153
rect 1003 85 1061 119
rect 1003 51 1015 85
rect 1049 51 1061 85
rect 1003 17 1061 51
rect 1003 -17 1015 17
rect 1049 -17 1061 17
rect 1003 -51 1061 -17
rect 1003 -85 1015 -51
rect 1049 -85 1061 -51
rect 1003 -119 1061 -85
rect 1003 -153 1015 -119
rect 1049 -153 1061 -119
rect 1003 -187 1061 -153
rect 1003 -221 1015 -187
rect 1049 -221 1061 -187
rect 1003 -255 1061 -221
rect 1003 -289 1015 -255
rect 1049 -289 1061 -255
rect 1003 -323 1061 -289
rect 1003 -357 1015 -323
rect 1049 -357 1061 -323
rect 1003 -391 1061 -357
rect 1003 -425 1015 -391
rect 1049 -425 1061 -391
rect 1003 -459 1061 -425
rect 1003 -493 1015 -459
rect 1049 -493 1061 -459
rect 1003 -527 1061 -493
rect 1003 -561 1015 -527
rect 1049 -561 1061 -527
rect 1003 -595 1061 -561
rect 1003 -629 1015 -595
rect 1049 -629 1061 -595
rect 1003 -663 1061 -629
rect 1003 -697 1015 -663
rect 1049 -697 1061 -663
rect 1003 -731 1061 -697
rect 1003 -765 1015 -731
rect 1049 -765 1061 -731
rect 1003 -800 1061 -765
rect 1261 765 1319 800
rect 1261 731 1273 765
rect 1307 731 1319 765
rect 1261 697 1319 731
rect 1261 663 1273 697
rect 1307 663 1319 697
rect 1261 629 1319 663
rect 1261 595 1273 629
rect 1307 595 1319 629
rect 1261 561 1319 595
rect 1261 527 1273 561
rect 1307 527 1319 561
rect 1261 493 1319 527
rect 1261 459 1273 493
rect 1307 459 1319 493
rect 1261 425 1319 459
rect 1261 391 1273 425
rect 1307 391 1319 425
rect 1261 357 1319 391
rect 1261 323 1273 357
rect 1307 323 1319 357
rect 1261 289 1319 323
rect 1261 255 1273 289
rect 1307 255 1319 289
rect 1261 221 1319 255
rect 1261 187 1273 221
rect 1307 187 1319 221
rect 1261 153 1319 187
rect 1261 119 1273 153
rect 1307 119 1319 153
rect 1261 85 1319 119
rect 1261 51 1273 85
rect 1307 51 1319 85
rect 1261 17 1319 51
rect 1261 -17 1273 17
rect 1307 -17 1319 17
rect 1261 -51 1319 -17
rect 1261 -85 1273 -51
rect 1307 -85 1319 -51
rect 1261 -119 1319 -85
rect 1261 -153 1273 -119
rect 1307 -153 1319 -119
rect 1261 -187 1319 -153
rect 1261 -221 1273 -187
rect 1307 -221 1319 -187
rect 1261 -255 1319 -221
rect 1261 -289 1273 -255
rect 1307 -289 1319 -255
rect 1261 -323 1319 -289
rect 1261 -357 1273 -323
rect 1307 -357 1319 -323
rect 1261 -391 1319 -357
rect 1261 -425 1273 -391
rect 1307 -425 1319 -391
rect 1261 -459 1319 -425
rect 1261 -493 1273 -459
rect 1307 -493 1319 -459
rect 1261 -527 1319 -493
rect 1261 -561 1273 -527
rect 1307 -561 1319 -527
rect 1261 -595 1319 -561
rect 1261 -629 1273 -595
rect 1307 -629 1319 -595
rect 1261 -663 1319 -629
rect 1261 -697 1273 -663
rect 1307 -697 1319 -663
rect 1261 -731 1319 -697
rect 1261 -765 1273 -731
rect 1307 -765 1319 -731
rect 1261 -800 1319 -765
<< pdiffc >>
rect -1307 731 -1273 765
rect -1307 663 -1273 697
rect -1307 595 -1273 629
rect -1307 527 -1273 561
rect -1307 459 -1273 493
rect -1307 391 -1273 425
rect -1307 323 -1273 357
rect -1307 255 -1273 289
rect -1307 187 -1273 221
rect -1307 119 -1273 153
rect -1307 51 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -51
rect -1307 -153 -1273 -119
rect -1307 -221 -1273 -187
rect -1307 -289 -1273 -255
rect -1307 -357 -1273 -323
rect -1307 -425 -1273 -391
rect -1307 -493 -1273 -459
rect -1307 -561 -1273 -527
rect -1307 -629 -1273 -595
rect -1307 -697 -1273 -663
rect -1307 -765 -1273 -731
rect -1049 731 -1015 765
rect -1049 663 -1015 697
rect -1049 595 -1015 629
rect -1049 527 -1015 561
rect -1049 459 -1015 493
rect -1049 391 -1015 425
rect -1049 323 -1015 357
rect -1049 255 -1015 289
rect -1049 187 -1015 221
rect -1049 119 -1015 153
rect -1049 51 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -51
rect -1049 -153 -1015 -119
rect -1049 -221 -1015 -187
rect -1049 -289 -1015 -255
rect -1049 -357 -1015 -323
rect -1049 -425 -1015 -391
rect -1049 -493 -1015 -459
rect -1049 -561 -1015 -527
rect -1049 -629 -1015 -595
rect -1049 -697 -1015 -663
rect -1049 -765 -1015 -731
rect -791 731 -757 765
rect -791 663 -757 697
rect -791 595 -757 629
rect -791 527 -757 561
rect -791 459 -757 493
rect -791 391 -757 425
rect -791 323 -757 357
rect -791 255 -757 289
rect -791 187 -757 221
rect -791 119 -757 153
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -791 -153 -757 -119
rect -791 -221 -757 -187
rect -791 -289 -757 -255
rect -791 -357 -757 -323
rect -791 -425 -757 -391
rect -791 -493 -757 -459
rect -791 -561 -757 -527
rect -791 -629 -757 -595
rect -791 -697 -757 -663
rect -791 -765 -757 -731
rect -533 731 -499 765
rect -533 663 -499 697
rect -533 595 -499 629
rect -533 527 -499 561
rect -533 459 -499 493
rect -533 391 -499 425
rect -533 323 -499 357
rect -533 255 -499 289
rect -533 187 -499 221
rect -533 119 -499 153
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -533 -153 -499 -119
rect -533 -221 -499 -187
rect -533 -289 -499 -255
rect -533 -357 -499 -323
rect -533 -425 -499 -391
rect -533 -493 -499 -459
rect -533 -561 -499 -527
rect -533 -629 -499 -595
rect -533 -697 -499 -663
rect -533 -765 -499 -731
rect -275 731 -241 765
rect -275 663 -241 697
rect -275 595 -241 629
rect -275 527 -241 561
rect -275 459 -241 493
rect -275 391 -241 425
rect -275 323 -241 357
rect -275 255 -241 289
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -275 -289 -241 -255
rect -275 -357 -241 -323
rect -275 -425 -241 -391
rect -275 -493 -241 -459
rect -275 -561 -241 -527
rect -275 -629 -241 -595
rect -275 -697 -241 -663
rect -275 -765 -241 -731
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect 241 731 275 765
rect 241 663 275 697
rect 241 595 275 629
rect 241 527 275 561
rect 241 459 275 493
rect 241 391 275 425
rect 241 323 275 357
rect 241 255 275 289
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect 241 -289 275 -255
rect 241 -357 275 -323
rect 241 -425 275 -391
rect 241 -493 275 -459
rect 241 -561 275 -527
rect 241 -629 275 -595
rect 241 -697 275 -663
rect 241 -765 275 -731
rect 499 731 533 765
rect 499 663 533 697
rect 499 595 533 629
rect 499 527 533 561
rect 499 459 533 493
rect 499 391 533 425
rect 499 323 533 357
rect 499 255 533 289
rect 499 187 533 221
rect 499 119 533 153
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 499 -153 533 -119
rect 499 -221 533 -187
rect 499 -289 533 -255
rect 499 -357 533 -323
rect 499 -425 533 -391
rect 499 -493 533 -459
rect 499 -561 533 -527
rect 499 -629 533 -595
rect 499 -697 533 -663
rect 499 -765 533 -731
rect 757 731 791 765
rect 757 663 791 697
rect 757 595 791 629
rect 757 527 791 561
rect 757 459 791 493
rect 757 391 791 425
rect 757 323 791 357
rect 757 255 791 289
rect 757 187 791 221
rect 757 119 791 153
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
rect 757 -153 791 -119
rect 757 -221 791 -187
rect 757 -289 791 -255
rect 757 -357 791 -323
rect 757 -425 791 -391
rect 757 -493 791 -459
rect 757 -561 791 -527
rect 757 -629 791 -595
rect 757 -697 791 -663
rect 757 -765 791 -731
rect 1015 731 1049 765
rect 1015 663 1049 697
rect 1015 595 1049 629
rect 1015 527 1049 561
rect 1015 459 1049 493
rect 1015 391 1049 425
rect 1015 323 1049 357
rect 1015 255 1049 289
rect 1015 187 1049 221
rect 1015 119 1049 153
rect 1015 51 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -51
rect 1015 -153 1049 -119
rect 1015 -221 1049 -187
rect 1015 -289 1049 -255
rect 1015 -357 1049 -323
rect 1015 -425 1049 -391
rect 1015 -493 1049 -459
rect 1015 -561 1049 -527
rect 1015 -629 1049 -595
rect 1015 -697 1049 -663
rect 1015 -765 1049 -731
rect 1273 731 1307 765
rect 1273 663 1307 697
rect 1273 595 1307 629
rect 1273 527 1307 561
rect 1273 459 1307 493
rect 1273 391 1307 425
rect 1273 323 1307 357
rect 1273 255 1307 289
rect 1273 187 1307 221
rect 1273 119 1307 153
rect 1273 51 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -51
rect 1273 -153 1307 -119
rect 1273 -221 1307 -187
rect 1273 -289 1307 -255
rect 1273 -357 1307 -323
rect 1273 -425 1307 -391
rect 1273 -493 1307 -459
rect 1273 -561 1307 -527
rect 1273 -629 1307 -595
rect 1273 -697 1307 -663
rect 1273 -765 1307 -731
<< nsubdiff >>
rect -1421 949 -1309 983
rect -1275 949 -1241 983
rect -1207 949 -1173 983
rect -1139 949 -1105 983
rect -1071 949 -1037 983
rect -1003 949 -969 983
rect -935 949 -901 983
rect -867 949 -833 983
rect -799 949 -765 983
rect -731 949 -697 983
rect -663 949 -629 983
rect -595 949 -561 983
rect -527 949 -493 983
rect -459 949 -425 983
rect -391 949 -357 983
rect -323 949 -289 983
rect -255 949 -221 983
rect -187 949 -153 983
rect -119 949 -85 983
rect -51 949 -17 983
rect 17 949 51 983
rect 85 949 119 983
rect 153 949 187 983
rect 221 949 255 983
rect 289 949 323 983
rect 357 949 391 983
rect 425 949 459 983
rect 493 949 527 983
rect 561 949 595 983
rect 629 949 663 983
rect 697 949 731 983
rect 765 949 799 983
rect 833 949 867 983
rect 901 949 935 983
rect 969 949 1003 983
rect 1037 949 1071 983
rect 1105 949 1139 983
rect 1173 949 1207 983
rect 1241 949 1275 983
rect 1309 949 1421 983
rect -1421 867 -1387 949
rect -1421 799 -1387 833
rect 1387 867 1421 949
rect -1421 731 -1387 765
rect -1421 663 -1387 697
rect -1421 595 -1387 629
rect -1421 527 -1387 561
rect -1421 459 -1387 493
rect -1421 391 -1387 425
rect -1421 323 -1387 357
rect -1421 255 -1387 289
rect -1421 187 -1387 221
rect -1421 119 -1387 153
rect -1421 51 -1387 85
rect -1421 -17 -1387 17
rect -1421 -85 -1387 -51
rect -1421 -153 -1387 -119
rect -1421 -221 -1387 -187
rect -1421 -289 -1387 -255
rect -1421 -357 -1387 -323
rect -1421 -425 -1387 -391
rect -1421 -493 -1387 -459
rect -1421 -561 -1387 -527
rect -1421 -629 -1387 -595
rect -1421 -697 -1387 -663
rect -1421 -765 -1387 -731
rect -1421 -833 -1387 -799
rect 1387 799 1421 833
rect 1387 731 1421 765
rect 1387 663 1421 697
rect 1387 595 1421 629
rect 1387 527 1421 561
rect 1387 459 1421 493
rect 1387 391 1421 425
rect 1387 323 1421 357
rect 1387 255 1421 289
rect 1387 187 1421 221
rect 1387 119 1421 153
rect 1387 51 1421 85
rect 1387 -17 1421 17
rect 1387 -85 1421 -51
rect 1387 -153 1421 -119
rect 1387 -221 1421 -187
rect 1387 -289 1421 -255
rect 1387 -357 1421 -323
rect 1387 -425 1421 -391
rect 1387 -493 1421 -459
rect 1387 -561 1421 -527
rect 1387 -629 1421 -595
rect 1387 -697 1421 -663
rect 1387 -765 1421 -731
rect -1421 -949 -1387 -867
rect 1387 -833 1421 -799
rect 1387 -949 1421 -867
rect -1421 -983 -1309 -949
rect -1275 -983 -1241 -949
rect -1207 -983 -1173 -949
rect -1139 -983 -1105 -949
rect -1071 -983 -1037 -949
rect -1003 -983 -969 -949
rect -935 -983 -901 -949
rect -867 -983 -833 -949
rect -799 -983 -765 -949
rect -731 -983 -697 -949
rect -663 -983 -629 -949
rect -595 -983 -561 -949
rect -527 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 527 -949
rect 561 -983 595 -949
rect 629 -983 663 -949
rect 697 -983 731 -949
rect 765 -983 799 -949
rect 833 -983 867 -949
rect 901 -983 935 -949
rect 969 -983 1003 -949
rect 1037 -983 1071 -949
rect 1105 -983 1139 -949
rect 1173 -983 1207 -949
rect 1241 -983 1275 -949
rect 1309 -983 1421 -949
<< nsubdiffcont >>
rect -1309 949 -1275 983
rect -1241 949 -1207 983
rect -1173 949 -1139 983
rect -1105 949 -1071 983
rect -1037 949 -1003 983
rect -969 949 -935 983
rect -901 949 -867 983
rect -833 949 -799 983
rect -765 949 -731 983
rect -697 949 -663 983
rect -629 949 -595 983
rect -561 949 -527 983
rect -493 949 -459 983
rect -425 949 -391 983
rect -357 949 -323 983
rect -289 949 -255 983
rect -221 949 -187 983
rect -153 949 -119 983
rect -85 949 -51 983
rect -17 949 17 983
rect 51 949 85 983
rect 119 949 153 983
rect 187 949 221 983
rect 255 949 289 983
rect 323 949 357 983
rect 391 949 425 983
rect 459 949 493 983
rect 527 949 561 983
rect 595 949 629 983
rect 663 949 697 983
rect 731 949 765 983
rect 799 949 833 983
rect 867 949 901 983
rect 935 949 969 983
rect 1003 949 1037 983
rect 1071 949 1105 983
rect 1139 949 1173 983
rect 1207 949 1241 983
rect 1275 949 1309 983
rect -1421 833 -1387 867
rect 1387 833 1421 867
rect -1421 765 -1387 799
rect -1421 697 -1387 731
rect -1421 629 -1387 663
rect -1421 561 -1387 595
rect -1421 493 -1387 527
rect -1421 425 -1387 459
rect -1421 357 -1387 391
rect -1421 289 -1387 323
rect -1421 221 -1387 255
rect -1421 153 -1387 187
rect -1421 85 -1387 119
rect -1421 17 -1387 51
rect -1421 -51 -1387 -17
rect -1421 -119 -1387 -85
rect -1421 -187 -1387 -153
rect -1421 -255 -1387 -221
rect -1421 -323 -1387 -289
rect -1421 -391 -1387 -357
rect -1421 -459 -1387 -425
rect -1421 -527 -1387 -493
rect -1421 -595 -1387 -561
rect -1421 -663 -1387 -629
rect -1421 -731 -1387 -697
rect -1421 -799 -1387 -765
rect 1387 765 1421 799
rect 1387 697 1421 731
rect 1387 629 1421 663
rect 1387 561 1421 595
rect 1387 493 1421 527
rect 1387 425 1421 459
rect 1387 357 1421 391
rect 1387 289 1421 323
rect 1387 221 1421 255
rect 1387 153 1421 187
rect 1387 85 1421 119
rect 1387 17 1421 51
rect 1387 -51 1421 -17
rect 1387 -119 1421 -85
rect 1387 -187 1421 -153
rect 1387 -255 1421 -221
rect 1387 -323 1421 -289
rect 1387 -391 1421 -357
rect 1387 -459 1421 -425
rect 1387 -527 1421 -493
rect 1387 -595 1421 -561
rect 1387 -663 1421 -629
rect 1387 -731 1421 -697
rect 1387 -799 1421 -765
rect -1421 -867 -1387 -833
rect 1387 -867 1421 -833
rect -1309 -983 -1275 -949
rect -1241 -983 -1207 -949
rect -1173 -983 -1139 -949
rect -1105 -983 -1071 -949
rect -1037 -983 -1003 -949
rect -969 -983 -935 -949
rect -901 -983 -867 -949
rect -833 -983 -799 -949
rect -765 -983 -731 -949
rect -697 -983 -663 -949
rect -629 -983 -595 -949
rect -561 -983 -527 -949
rect -493 -983 -459 -949
rect -425 -983 -391 -949
rect -357 -983 -323 -949
rect -289 -983 -255 -949
rect -221 -983 -187 -949
rect -153 -983 -119 -949
rect -85 -983 -51 -949
rect -17 -983 17 -949
rect 51 -983 85 -949
rect 119 -983 153 -949
rect 187 -983 221 -949
rect 255 -983 289 -949
rect 323 -983 357 -949
rect 391 -983 425 -949
rect 459 -983 493 -949
rect 527 -983 561 -949
rect 595 -983 629 -949
rect 663 -983 697 -949
rect 731 -983 765 -949
rect 799 -983 833 -949
rect 867 -983 901 -949
rect 935 -983 969 -949
rect 1003 -983 1037 -949
rect 1071 -983 1105 -949
rect 1139 -983 1173 -949
rect 1207 -983 1241 -949
rect 1275 -983 1309 -949
<< poly >>
rect -1261 881 -1061 897
rect -1261 847 -1212 881
rect -1178 847 -1144 881
rect -1110 847 -1061 881
rect -1261 800 -1061 847
rect -1003 881 -803 897
rect -1003 847 -954 881
rect -920 847 -886 881
rect -852 847 -803 881
rect -1003 800 -803 847
rect -745 881 -545 897
rect -745 847 -696 881
rect -662 847 -628 881
rect -594 847 -545 881
rect -745 800 -545 847
rect -487 881 -287 897
rect -487 847 -438 881
rect -404 847 -370 881
rect -336 847 -287 881
rect -487 800 -287 847
rect -229 881 -29 897
rect -229 847 -180 881
rect -146 847 -112 881
rect -78 847 -29 881
rect -229 800 -29 847
rect 29 881 229 897
rect 29 847 78 881
rect 112 847 146 881
rect 180 847 229 881
rect 29 800 229 847
rect 287 881 487 897
rect 287 847 336 881
rect 370 847 404 881
rect 438 847 487 881
rect 287 800 487 847
rect 545 881 745 897
rect 545 847 594 881
rect 628 847 662 881
rect 696 847 745 881
rect 545 800 745 847
rect 803 881 1003 897
rect 803 847 852 881
rect 886 847 920 881
rect 954 847 1003 881
rect 803 800 1003 847
rect 1061 881 1261 897
rect 1061 847 1110 881
rect 1144 847 1178 881
rect 1212 847 1261 881
rect 1061 800 1261 847
rect -1261 -847 -1061 -800
rect -1261 -881 -1212 -847
rect -1178 -881 -1144 -847
rect -1110 -881 -1061 -847
rect -1261 -897 -1061 -881
rect -1003 -847 -803 -800
rect -1003 -881 -954 -847
rect -920 -881 -886 -847
rect -852 -881 -803 -847
rect -1003 -897 -803 -881
rect -745 -847 -545 -800
rect -745 -881 -696 -847
rect -662 -881 -628 -847
rect -594 -881 -545 -847
rect -745 -897 -545 -881
rect -487 -847 -287 -800
rect -487 -881 -438 -847
rect -404 -881 -370 -847
rect -336 -881 -287 -847
rect -487 -897 -287 -881
rect -229 -847 -29 -800
rect -229 -881 -180 -847
rect -146 -881 -112 -847
rect -78 -881 -29 -847
rect -229 -897 -29 -881
rect 29 -847 229 -800
rect 29 -881 78 -847
rect 112 -881 146 -847
rect 180 -881 229 -847
rect 29 -897 229 -881
rect 287 -847 487 -800
rect 287 -881 336 -847
rect 370 -881 404 -847
rect 438 -881 487 -847
rect 287 -897 487 -881
rect 545 -847 745 -800
rect 545 -881 594 -847
rect 628 -881 662 -847
rect 696 -881 745 -847
rect 545 -897 745 -881
rect 803 -847 1003 -800
rect 803 -881 852 -847
rect 886 -881 920 -847
rect 954 -881 1003 -847
rect 803 -897 1003 -881
rect 1061 -847 1261 -800
rect 1061 -881 1110 -847
rect 1144 -881 1178 -847
rect 1212 -881 1261 -847
rect 1061 -897 1261 -881
<< polycont >>
rect -1212 847 -1178 881
rect -1144 847 -1110 881
rect -954 847 -920 881
rect -886 847 -852 881
rect -696 847 -662 881
rect -628 847 -594 881
rect -438 847 -404 881
rect -370 847 -336 881
rect -180 847 -146 881
rect -112 847 -78 881
rect 78 847 112 881
rect 146 847 180 881
rect 336 847 370 881
rect 404 847 438 881
rect 594 847 628 881
rect 662 847 696 881
rect 852 847 886 881
rect 920 847 954 881
rect 1110 847 1144 881
rect 1178 847 1212 881
rect -1212 -881 -1178 -847
rect -1144 -881 -1110 -847
rect -954 -881 -920 -847
rect -886 -881 -852 -847
rect -696 -881 -662 -847
rect -628 -881 -594 -847
rect -438 -881 -404 -847
rect -370 -881 -336 -847
rect -180 -881 -146 -847
rect -112 -881 -78 -847
rect 78 -881 112 -847
rect 146 -881 180 -847
rect 336 -881 370 -847
rect 404 -881 438 -847
rect 594 -881 628 -847
rect 662 -881 696 -847
rect 852 -881 886 -847
rect 920 -881 954 -847
rect 1110 -881 1144 -847
rect 1178 -881 1212 -847
<< locali >>
rect -1421 949 -1309 983
rect -1275 949 -1241 983
rect -1207 949 -1173 983
rect -1139 949 -1105 983
rect -1071 949 -1037 983
rect -1003 949 -969 983
rect -935 949 -901 983
rect -867 949 -833 983
rect -799 949 -765 983
rect -731 949 -697 983
rect -663 949 -629 983
rect -595 949 -561 983
rect -527 949 -493 983
rect -459 949 -425 983
rect -391 949 -357 983
rect -323 949 -289 983
rect -255 949 -221 983
rect -187 949 -153 983
rect -119 949 -85 983
rect -51 949 -17 983
rect 17 949 51 983
rect 85 949 119 983
rect 153 949 187 983
rect 221 949 255 983
rect 289 949 323 983
rect 357 949 391 983
rect 425 949 459 983
rect 493 949 527 983
rect 561 949 595 983
rect 629 949 663 983
rect 697 949 731 983
rect 765 949 799 983
rect 833 949 867 983
rect 901 949 935 983
rect 969 949 1003 983
rect 1037 949 1071 983
rect 1105 949 1139 983
rect 1173 949 1207 983
rect 1241 949 1275 983
rect 1309 949 1421 983
rect -1421 867 -1387 949
rect -1261 847 -1214 881
rect -1178 847 -1144 881
rect -1108 847 -1061 881
rect -1003 847 -956 881
rect -920 847 -886 881
rect -850 847 -803 881
rect -745 847 -698 881
rect -662 847 -628 881
rect -592 847 -545 881
rect -487 847 -440 881
rect -404 847 -370 881
rect -334 847 -287 881
rect -229 847 -182 881
rect -146 847 -112 881
rect -76 847 -29 881
rect 29 847 76 881
rect 112 847 146 881
rect 182 847 229 881
rect 287 847 334 881
rect 370 847 404 881
rect 440 847 487 881
rect 545 847 592 881
rect 628 847 662 881
rect 698 847 745 881
rect 803 847 850 881
rect 886 847 920 881
rect 956 847 1003 881
rect 1061 847 1108 881
rect 1144 847 1178 881
rect 1214 847 1261 881
rect 1387 867 1421 949
rect -1421 799 -1387 833
rect -1421 731 -1387 765
rect -1421 663 -1387 697
rect -1421 595 -1387 629
rect -1421 527 -1387 561
rect -1421 459 -1387 493
rect -1421 391 -1387 425
rect -1421 323 -1387 357
rect -1421 255 -1387 289
rect -1421 187 -1387 221
rect -1421 119 -1387 153
rect -1421 51 -1387 85
rect -1421 -17 -1387 17
rect -1421 -85 -1387 -51
rect -1421 -153 -1387 -119
rect -1421 -221 -1387 -187
rect -1421 -289 -1387 -255
rect -1421 -357 -1387 -323
rect -1421 -425 -1387 -391
rect -1421 -493 -1387 -459
rect -1421 -561 -1387 -527
rect -1421 -629 -1387 -595
rect -1421 -697 -1387 -663
rect -1421 -765 -1387 -731
rect -1421 -833 -1387 -799
rect -1307 773 -1273 804
rect -1307 701 -1273 731
rect -1307 629 -1273 663
rect -1307 561 -1273 595
rect -1307 493 -1273 523
rect -1307 425 -1273 451
rect -1307 357 -1273 379
rect -1307 289 -1273 307
rect -1307 221 -1273 235
rect -1307 153 -1273 163
rect -1307 85 -1273 91
rect -1307 17 -1273 19
rect -1307 -19 -1273 -17
rect -1307 -91 -1273 -85
rect -1307 -163 -1273 -153
rect -1307 -235 -1273 -221
rect -1307 -307 -1273 -289
rect -1307 -379 -1273 -357
rect -1307 -451 -1273 -425
rect -1307 -523 -1273 -493
rect -1307 -595 -1273 -561
rect -1307 -663 -1273 -629
rect -1307 -731 -1273 -701
rect -1307 -804 -1273 -773
rect -1049 773 -1015 804
rect -1049 701 -1015 731
rect -1049 629 -1015 663
rect -1049 561 -1015 595
rect -1049 493 -1015 523
rect -1049 425 -1015 451
rect -1049 357 -1015 379
rect -1049 289 -1015 307
rect -1049 221 -1015 235
rect -1049 153 -1015 163
rect -1049 85 -1015 91
rect -1049 17 -1015 19
rect -1049 -19 -1015 -17
rect -1049 -91 -1015 -85
rect -1049 -163 -1015 -153
rect -1049 -235 -1015 -221
rect -1049 -307 -1015 -289
rect -1049 -379 -1015 -357
rect -1049 -451 -1015 -425
rect -1049 -523 -1015 -493
rect -1049 -595 -1015 -561
rect -1049 -663 -1015 -629
rect -1049 -731 -1015 -701
rect -1049 -804 -1015 -773
rect -791 773 -757 804
rect -791 701 -757 731
rect -791 629 -757 663
rect -791 561 -757 595
rect -791 493 -757 523
rect -791 425 -757 451
rect -791 357 -757 379
rect -791 289 -757 307
rect -791 221 -757 235
rect -791 153 -757 163
rect -791 85 -757 91
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -91 -757 -85
rect -791 -163 -757 -153
rect -791 -235 -757 -221
rect -791 -307 -757 -289
rect -791 -379 -757 -357
rect -791 -451 -757 -425
rect -791 -523 -757 -493
rect -791 -595 -757 -561
rect -791 -663 -757 -629
rect -791 -731 -757 -701
rect -791 -804 -757 -773
rect -533 773 -499 804
rect -533 701 -499 731
rect -533 629 -499 663
rect -533 561 -499 595
rect -533 493 -499 523
rect -533 425 -499 451
rect -533 357 -499 379
rect -533 289 -499 307
rect -533 221 -499 235
rect -533 153 -499 163
rect -533 85 -499 91
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -91 -499 -85
rect -533 -163 -499 -153
rect -533 -235 -499 -221
rect -533 -307 -499 -289
rect -533 -379 -499 -357
rect -533 -451 -499 -425
rect -533 -523 -499 -493
rect -533 -595 -499 -561
rect -533 -663 -499 -629
rect -533 -731 -499 -701
rect -533 -804 -499 -773
rect -275 773 -241 804
rect -275 701 -241 731
rect -275 629 -241 663
rect -275 561 -241 595
rect -275 493 -241 523
rect -275 425 -241 451
rect -275 357 -241 379
rect -275 289 -241 307
rect -275 221 -241 235
rect -275 153 -241 163
rect -275 85 -241 91
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -91 -241 -85
rect -275 -163 -241 -153
rect -275 -235 -241 -221
rect -275 -307 -241 -289
rect -275 -379 -241 -357
rect -275 -451 -241 -425
rect -275 -523 -241 -493
rect -275 -595 -241 -561
rect -275 -663 -241 -629
rect -275 -731 -241 -701
rect -275 -804 -241 -773
rect -17 773 17 804
rect -17 701 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -701
rect -17 -804 17 -773
rect 241 773 275 804
rect 241 701 275 731
rect 241 629 275 663
rect 241 561 275 595
rect 241 493 275 523
rect 241 425 275 451
rect 241 357 275 379
rect 241 289 275 307
rect 241 221 275 235
rect 241 153 275 163
rect 241 85 275 91
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -91 275 -85
rect 241 -163 275 -153
rect 241 -235 275 -221
rect 241 -307 275 -289
rect 241 -379 275 -357
rect 241 -451 275 -425
rect 241 -523 275 -493
rect 241 -595 275 -561
rect 241 -663 275 -629
rect 241 -731 275 -701
rect 241 -804 275 -773
rect 499 773 533 804
rect 499 701 533 731
rect 499 629 533 663
rect 499 561 533 595
rect 499 493 533 523
rect 499 425 533 451
rect 499 357 533 379
rect 499 289 533 307
rect 499 221 533 235
rect 499 153 533 163
rect 499 85 533 91
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -91 533 -85
rect 499 -163 533 -153
rect 499 -235 533 -221
rect 499 -307 533 -289
rect 499 -379 533 -357
rect 499 -451 533 -425
rect 499 -523 533 -493
rect 499 -595 533 -561
rect 499 -663 533 -629
rect 499 -731 533 -701
rect 499 -804 533 -773
rect 757 773 791 804
rect 757 701 791 731
rect 757 629 791 663
rect 757 561 791 595
rect 757 493 791 523
rect 757 425 791 451
rect 757 357 791 379
rect 757 289 791 307
rect 757 221 791 235
rect 757 153 791 163
rect 757 85 791 91
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -91 791 -85
rect 757 -163 791 -153
rect 757 -235 791 -221
rect 757 -307 791 -289
rect 757 -379 791 -357
rect 757 -451 791 -425
rect 757 -523 791 -493
rect 757 -595 791 -561
rect 757 -663 791 -629
rect 757 -731 791 -701
rect 757 -804 791 -773
rect 1015 773 1049 804
rect 1015 701 1049 731
rect 1015 629 1049 663
rect 1015 561 1049 595
rect 1015 493 1049 523
rect 1015 425 1049 451
rect 1015 357 1049 379
rect 1015 289 1049 307
rect 1015 221 1049 235
rect 1015 153 1049 163
rect 1015 85 1049 91
rect 1015 17 1049 19
rect 1015 -19 1049 -17
rect 1015 -91 1049 -85
rect 1015 -163 1049 -153
rect 1015 -235 1049 -221
rect 1015 -307 1049 -289
rect 1015 -379 1049 -357
rect 1015 -451 1049 -425
rect 1015 -523 1049 -493
rect 1015 -595 1049 -561
rect 1015 -663 1049 -629
rect 1015 -731 1049 -701
rect 1015 -804 1049 -773
rect 1273 773 1307 804
rect 1273 701 1307 731
rect 1273 629 1307 663
rect 1273 561 1307 595
rect 1273 493 1307 523
rect 1273 425 1307 451
rect 1273 357 1307 379
rect 1273 289 1307 307
rect 1273 221 1307 235
rect 1273 153 1307 163
rect 1273 85 1307 91
rect 1273 17 1307 19
rect 1273 -19 1307 -17
rect 1273 -91 1307 -85
rect 1273 -163 1307 -153
rect 1273 -235 1307 -221
rect 1273 -307 1307 -289
rect 1273 -379 1307 -357
rect 1273 -451 1307 -425
rect 1273 -523 1307 -493
rect 1273 -595 1307 -561
rect 1273 -663 1307 -629
rect 1273 -731 1307 -701
rect 1273 -804 1307 -773
rect 1387 799 1421 833
rect 1387 731 1421 765
rect 1387 663 1421 697
rect 1387 595 1421 629
rect 1387 527 1421 561
rect 1387 459 1421 493
rect 1387 391 1421 425
rect 1387 323 1421 357
rect 1387 255 1421 289
rect 1387 187 1421 221
rect 1387 119 1421 153
rect 1387 51 1421 85
rect 1387 -17 1421 17
rect 1387 -85 1421 -51
rect 1387 -153 1421 -119
rect 1387 -221 1421 -187
rect 1387 -289 1421 -255
rect 1387 -357 1421 -323
rect 1387 -425 1421 -391
rect 1387 -493 1421 -459
rect 1387 -561 1421 -527
rect 1387 -629 1421 -595
rect 1387 -697 1421 -663
rect 1387 -765 1421 -731
rect 1387 -833 1421 -799
rect -1421 -949 -1387 -867
rect -1261 -881 -1214 -847
rect -1178 -881 -1144 -847
rect -1108 -881 -1061 -847
rect -1003 -881 -956 -847
rect -920 -881 -886 -847
rect -850 -881 -803 -847
rect -745 -881 -698 -847
rect -662 -881 -628 -847
rect -592 -881 -545 -847
rect -487 -881 -440 -847
rect -404 -881 -370 -847
rect -334 -881 -287 -847
rect -229 -881 -182 -847
rect -146 -881 -112 -847
rect -76 -881 -29 -847
rect 29 -881 76 -847
rect 112 -881 146 -847
rect 182 -881 229 -847
rect 287 -881 334 -847
rect 370 -881 404 -847
rect 440 -881 487 -847
rect 545 -881 592 -847
rect 628 -881 662 -847
rect 698 -881 745 -847
rect 803 -881 850 -847
rect 886 -881 920 -847
rect 956 -881 1003 -847
rect 1061 -881 1108 -847
rect 1144 -881 1178 -847
rect 1214 -881 1261 -847
rect 1387 -949 1421 -867
rect -1421 -983 -1309 -949
rect -1275 -983 -1241 -949
rect -1207 -983 -1173 -949
rect -1139 -983 -1105 -949
rect -1071 -983 -1037 -949
rect -1003 -983 -969 -949
rect -935 -983 -901 -949
rect -867 -983 -833 -949
rect -799 -983 -765 -949
rect -731 -983 -697 -949
rect -663 -983 -629 -949
rect -595 -983 -561 -949
rect -527 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 527 -949
rect 561 -983 595 -949
rect 629 -983 663 -949
rect 697 -983 731 -949
rect 765 -983 799 -949
rect 833 -983 867 -949
rect 901 -983 935 -949
rect 969 -983 1003 -949
rect 1037 -983 1071 -949
rect 1105 -983 1139 -949
rect 1173 -983 1207 -949
rect 1241 -983 1275 -949
rect 1309 -983 1421 -949
<< viali >>
rect -1214 847 -1212 881
rect -1212 847 -1180 881
rect -1142 847 -1110 881
rect -1110 847 -1108 881
rect -956 847 -954 881
rect -954 847 -922 881
rect -884 847 -852 881
rect -852 847 -850 881
rect -698 847 -696 881
rect -696 847 -664 881
rect -626 847 -594 881
rect -594 847 -592 881
rect -440 847 -438 881
rect -438 847 -406 881
rect -368 847 -336 881
rect -336 847 -334 881
rect -182 847 -180 881
rect -180 847 -148 881
rect -110 847 -78 881
rect -78 847 -76 881
rect 76 847 78 881
rect 78 847 110 881
rect 148 847 180 881
rect 180 847 182 881
rect 334 847 336 881
rect 336 847 368 881
rect 406 847 438 881
rect 438 847 440 881
rect 592 847 594 881
rect 594 847 626 881
rect 664 847 696 881
rect 696 847 698 881
rect 850 847 852 881
rect 852 847 884 881
rect 922 847 954 881
rect 954 847 956 881
rect 1108 847 1110 881
rect 1110 847 1142 881
rect 1180 847 1212 881
rect 1212 847 1214 881
rect -1307 765 -1273 773
rect -1307 739 -1273 765
rect -1307 697 -1273 701
rect -1307 667 -1273 697
rect -1307 595 -1273 629
rect -1307 527 -1273 557
rect -1307 523 -1273 527
rect -1307 459 -1273 485
rect -1307 451 -1273 459
rect -1307 391 -1273 413
rect -1307 379 -1273 391
rect -1307 323 -1273 341
rect -1307 307 -1273 323
rect -1307 255 -1273 269
rect -1307 235 -1273 255
rect -1307 187 -1273 197
rect -1307 163 -1273 187
rect -1307 119 -1273 125
rect -1307 91 -1273 119
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1307 -119 -1273 -91
rect -1307 -125 -1273 -119
rect -1307 -187 -1273 -163
rect -1307 -197 -1273 -187
rect -1307 -255 -1273 -235
rect -1307 -269 -1273 -255
rect -1307 -323 -1273 -307
rect -1307 -341 -1273 -323
rect -1307 -391 -1273 -379
rect -1307 -413 -1273 -391
rect -1307 -459 -1273 -451
rect -1307 -485 -1273 -459
rect -1307 -527 -1273 -523
rect -1307 -557 -1273 -527
rect -1307 -629 -1273 -595
rect -1307 -697 -1273 -667
rect -1307 -701 -1273 -697
rect -1307 -765 -1273 -739
rect -1307 -773 -1273 -765
rect -1049 765 -1015 773
rect -1049 739 -1015 765
rect -1049 697 -1015 701
rect -1049 667 -1015 697
rect -1049 595 -1015 629
rect -1049 527 -1015 557
rect -1049 523 -1015 527
rect -1049 459 -1015 485
rect -1049 451 -1015 459
rect -1049 391 -1015 413
rect -1049 379 -1015 391
rect -1049 323 -1015 341
rect -1049 307 -1015 323
rect -1049 255 -1015 269
rect -1049 235 -1015 255
rect -1049 187 -1015 197
rect -1049 163 -1015 187
rect -1049 119 -1015 125
rect -1049 91 -1015 119
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -1049 -119 -1015 -91
rect -1049 -125 -1015 -119
rect -1049 -187 -1015 -163
rect -1049 -197 -1015 -187
rect -1049 -255 -1015 -235
rect -1049 -269 -1015 -255
rect -1049 -323 -1015 -307
rect -1049 -341 -1015 -323
rect -1049 -391 -1015 -379
rect -1049 -413 -1015 -391
rect -1049 -459 -1015 -451
rect -1049 -485 -1015 -459
rect -1049 -527 -1015 -523
rect -1049 -557 -1015 -527
rect -1049 -629 -1015 -595
rect -1049 -697 -1015 -667
rect -1049 -701 -1015 -697
rect -1049 -765 -1015 -739
rect -1049 -773 -1015 -765
rect -791 765 -757 773
rect -791 739 -757 765
rect -791 697 -757 701
rect -791 667 -757 697
rect -791 595 -757 629
rect -791 527 -757 557
rect -791 523 -757 527
rect -791 459 -757 485
rect -791 451 -757 459
rect -791 391 -757 413
rect -791 379 -757 391
rect -791 323 -757 341
rect -791 307 -757 323
rect -791 255 -757 269
rect -791 235 -757 255
rect -791 187 -757 197
rect -791 163 -757 187
rect -791 119 -757 125
rect -791 91 -757 119
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -791 -119 -757 -91
rect -791 -125 -757 -119
rect -791 -187 -757 -163
rect -791 -197 -757 -187
rect -791 -255 -757 -235
rect -791 -269 -757 -255
rect -791 -323 -757 -307
rect -791 -341 -757 -323
rect -791 -391 -757 -379
rect -791 -413 -757 -391
rect -791 -459 -757 -451
rect -791 -485 -757 -459
rect -791 -527 -757 -523
rect -791 -557 -757 -527
rect -791 -629 -757 -595
rect -791 -697 -757 -667
rect -791 -701 -757 -697
rect -791 -765 -757 -739
rect -791 -773 -757 -765
rect -533 765 -499 773
rect -533 739 -499 765
rect -533 697 -499 701
rect -533 667 -499 697
rect -533 595 -499 629
rect -533 527 -499 557
rect -533 523 -499 527
rect -533 459 -499 485
rect -533 451 -499 459
rect -533 391 -499 413
rect -533 379 -499 391
rect -533 323 -499 341
rect -533 307 -499 323
rect -533 255 -499 269
rect -533 235 -499 255
rect -533 187 -499 197
rect -533 163 -499 187
rect -533 119 -499 125
rect -533 91 -499 119
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -533 -119 -499 -91
rect -533 -125 -499 -119
rect -533 -187 -499 -163
rect -533 -197 -499 -187
rect -533 -255 -499 -235
rect -533 -269 -499 -255
rect -533 -323 -499 -307
rect -533 -341 -499 -323
rect -533 -391 -499 -379
rect -533 -413 -499 -391
rect -533 -459 -499 -451
rect -533 -485 -499 -459
rect -533 -527 -499 -523
rect -533 -557 -499 -527
rect -533 -629 -499 -595
rect -533 -697 -499 -667
rect -533 -701 -499 -697
rect -533 -765 -499 -739
rect -533 -773 -499 -765
rect -275 765 -241 773
rect -275 739 -241 765
rect -275 697 -241 701
rect -275 667 -241 697
rect -275 595 -241 629
rect -275 527 -241 557
rect -275 523 -241 527
rect -275 459 -241 485
rect -275 451 -241 459
rect -275 391 -241 413
rect -275 379 -241 391
rect -275 323 -241 341
rect -275 307 -241 323
rect -275 255 -241 269
rect -275 235 -241 255
rect -275 187 -241 197
rect -275 163 -241 187
rect -275 119 -241 125
rect -275 91 -241 119
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -275 -119 -241 -91
rect -275 -125 -241 -119
rect -275 -187 -241 -163
rect -275 -197 -241 -187
rect -275 -255 -241 -235
rect -275 -269 -241 -255
rect -275 -323 -241 -307
rect -275 -341 -241 -323
rect -275 -391 -241 -379
rect -275 -413 -241 -391
rect -275 -459 -241 -451
rect -275 -485 -241 -459
rect -275 -527 -241 -523
rect -275 -557 -241 -527
rect -275 -629 -241 -595
rect -275 -697 -241 -667
rect -275 -701 -241 -697
rect -275 -765 -241 -739
rect -275 -773 -241 -765
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect 241 765 275 773
rect 241 739 275 765
rect 241 697 275 701
rect 241 667 275 697
rect 241 595 275 629
rect 241 527 275 557
rect 241 523 275 527
rect 241 459 275 485
rect 241 451 275 459
rect 241 391 275 413
rect 241 379 275 391
rect 241 323 275 341
rect 241 307 275 323
rect 241 255 275 269
rect 241 235 275 255
rect 241 187 275 197
rect 241 163 275 187
rect 241 119 275 125
rect 241 91 275 119
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 241 -119 275 -91
rect 241 -125 275 -119
rect 241 -187 275 -163
rect 241 -197 275 -187
rect 241 -255 275 -235
rect 241 -269 275 -255
rect 241 -323 275 -307
rect 241 -341 275 -323
rect 241 -391 275 -379
rect 241 -413 275 -391
rect 241 -459 275 -451
rect 241 -485 275 -459
rect 241 -527 275 -523
rect 241 -557 275 -527
rect 241 -629 275 -595
rect 241 -697 275 -667
rect 241 -701 275 -697
rect 241 -765 275 -739
rect 241 -773 275 -765
rect 499 765 533 773
rect 499 739 533 765
rect 499 697 533 701
rect 499 667 533 697
rect 499 595 533 629
rect 499 527 533 557
rect 499 523 533 527
rect 499 459 533 485
rect 499 451 533 459
rect 499 391 533 413
rect 499 379 533 391
rect 499 323 533 341
rect 499 307 533 323
rect 499 255 533 269
rect 499 235 533 255
rect 499 187 533 197
rect 499 163 533 187
rect 499 119 533 125
rect 499 91 533 119
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 499 -119 533 -91
rect 499 -125 533 -119
rect 499 -187 533 -163
rect 499 -197 533 -187
rect 499 -255 533 -235
rect 499 -269 533 -255
rect 499 -323 533 -307
rect 499 -341 533 -323
rect 499 -391 533 -379
rect 499 -413 533 -391
rect 499 -459 533 -451
rect 499 -485 533 -459
rect 499 -527 533 -523
rect 499 -557 533 -527
rect 499 -629 533 -595
rect 499 -697 533 -667
rect 499 -701 533 -697
rect 499 -765 533 -739
rect 499 -773 533 -765
rect 757 765 791 773
rect 757 739 791 765
rect 757 697 791 701
rect 757 667 791 697
rect 757 595 791 629
rect 757 527 791 557
rect 757 523 791 527
rect 757 459 791 485
rect 757 451 791 459
rect 757 391 791 413
rect 757 379 791 391
rect 757 323 791 341
rect 757 307 791 323
rect 757 255 791 269
rect 757 235 791 255
rect 757 187 791 197
rect 757 163 791 187
rect 757 119 791 125
rect 757 91 791 119
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 757 -119 791 -91
rect 757 -125 791 -119
rect 757 -187 791 -163
rect 757 -197 791 -187
rect 757 -255 791 -235
rect 757 -269 791 -255
rect 757 -323 791 -307
rect 757 -341 791 -323
rect 757 -391 791 -379
rect 757 -413 791 -391
rect 757 -459 791 -451
rect 757 -485 791 -459
rect 757 -527 791 -523
rect 757 -557 791 -527
rect 757 -629 791 -595
rect 757 -697 791 -667
rect 757 -701 791 -697
rect 757 -765 791 -739
rect 757 -773 791 -765
rect 1015 765 1049 773
rect 1015 739 1049 765
rect 1015 697 1049 701
rect 1015 667 1049 697
rect 1015 595 1049 629
rect 1015 527 1049 557
rect 1015 523 1049 527
rect 1015 459 1049 485
rect 1015 451 1049 459
rect 1015 391 1049 413
rect 1015 379 1049 391
rect 1015 323 1049 341
rect 1015 307 1049 323
rect 1015 255 1049 269
rect 1015 235 1049 255
rect 1015 187 1049 197
rect 1015 163 1049 187
rect 1015 119 1049 125
rect 1015 91 1049 119
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1015 -119 1049 -91
rect 1015 -125 1049 -119
rect 1015 -187 1049 -163
rect 1015 -197 1049 -187
rect 1015 -255 1049 -235
rect 1015 -269 1049 -255
rect 1015 -323 1049 -307
rect 1015 -341 1049 -323
rect 1015 -391 1049 -379
rect 1015 -413 1049 -391
rect 1015 -459 1049 -451
rect 1015 -485 1049 -459
rect 1015 -527 1049 -523
rect 1015 -557 1049 -527
rect 1015 -629 1049 -595
rect 1015 -697 1049 -667
rect 1015 -701 1049 -697
rect 1015 -765 1049 -739
rect 1015 -773 1049 -765
rect 1273 765 1307 773
rect 1273 739 1307 765
rect 1273 697 1307 701
rect 1273 667 1307 697
rect 1273 595 1307 629
rect 1273 527 1307 557
rect 1273 523 1307 527
rect 1273 459 1307 485
rect 1273 451 1307 459
rect 1273 391 1307 413
rect 1273 379 1307 391
rect 1273 323 1307 341
rect 1273 307 1307 323
rect 1273 255 1307 269
rect 1273 235 1307 255
rect 1273 187 1307 197
rect 1273 163 1307 187
rect 1273 119 1307 125
rect 1273 91 1307 119
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect 1273 -119 1307 -91
rect 1273 -125 1307 -119
rect 1273 -187 1307 -163
rect 1273 -197 1307 -187
rect 1273 -255 1307 -235
rect 1273 -269 1307 -255
rect 1273 -323 1307 -307
rect 1273 -341 1307 -323
rect 1273 -391 1307 -379
rect 1273 -413 1307 -391
rect 1273 -459 1307 -451
rect 1273 -485 1307 -459
rect 1273 -527 1307 -523
rect 1273 -557 1307 -527
rect 1273 -629 1307 -595
rect 1273 -697 1307 -667
rect 1273 -701 1307 -697
rect 1273 -765 1307 -739
rect 1273 -773 1307 -765
rect -1214 -881 -1212 -847
rect -1212 -881 -1180 -847
rect -1142 -881 -1110 -847
rect -1110 -881 -1108 -847
rect -956 -881 -954 -847
rect -954 -881 -922 -847
rect -884 -881 -852 -847
rect -852 -881 -850 -847
rect -698 -881 -696 -847
rect -696 -881 -664 -847
rect -626 -881 -594 -847
rect -594 -881 -592 -847
rect -440 -881 -438 -847
rect -438 -881 -406 -847
rect -368 -881 -336 -847
rect -336 -881 -334 -847
rect -182 -881 -180 -847
rect -180 -881 -148 -847
rect -110 -881 -78 -847
rect -78 -881 -76 -847
rect 76 -881 78 -847
rect 78 -881 110 -847
rect 148 -881 180 -847
rect 180 -881 182 -847
rect 334 -881 336 -847
rect 336 -881 368 -847
rect 406 -881 438 -847
rect 438 -881 440 -847
rect 592 -881 594 -847
rect 594 -881 626 -847
rect 664 -881 696 -847
rect 696 -881 698 -847
rect 850 -881 852 -847
rect 852 -881 884 -847
rect 922 -881 954 -847
rect 954 -881 956 -847
rect 1108 -881 1110 -847
rect 1110 -881 1142 -847
rect 1180 -881 1212 -847
rect 1212 -881 1214 -847
<< metal1 >>
rect -1257 881 -1065 887
rect -1257 847 -1214 881
rect -1180 847 -1142 881
rect -1108 847 -1065 881
rect -1257 841 -1065 847
rect -999 881 -807 887
rect -999 847 -956 881
rect -922 847 -884 881
rect -850 847 -807 881
rect -999 841 -807 847
rect -741 881 -549 887
rect -741 847 -698 881
rect -664 847 -626 881
rect -592 847 -549 881
rect -741 841 -549 847
rect -483 881 -291 887
rect -483 847 -440 881
rect -406 847 -368 881
rect -334 847 -291 881
rect -483 841 -291 847
rect -225 881 -33 887
rect -225 847 -182 881
rect -148 847 -110 881
rect -76 847 -33 881
rect -225 841 -33 847
rect 33 881 225 887
rect 33 847 76 881
rect 110 847 148 881
rect 182 847 225 881
rect 33 841 225 847
rect 291 881 483 887
rect 291 847 334 881
rect 368 847 406 881
rect 440 847 483 881
rect 291 841 483 847
rect 549 881 741 887
rect 549 847 592 881
rect 626 847 664 881
rect 698 847 741 881
rect 549 841 741 847
rect 807 881 999 887
rect 807 847 850 881
rect 884 847 922 881
rect 956 847 999 881
rect 807 841 999 847
rect 1065 881 1257 887
rect 1065 847 1108 881
rect 1142 847 1180 881
rect 1214 847 1257 881
rect 1065 841 1257 847
rect -1313 773 -1267 800
rect -1313 739 -1307 773
rect -1273 739 -1267 773
rect -1313 701 -1267 739
rect -1313 667 -1307 701
rect -1273 667 -1267 701
rect -1313 629 -1267 667
rect -1313 595 -1307 629
rect -1273 595 -1267 629
rect -1313 557 -1267 595
rect -1313 523 -1307 557
rect -1273 523 -1267 557
rect -1313 485 -1267 523
rect -1313 451 -1307 485
rect -1273 451 -1267 485
rect -1313 413 -1267 451
rect -1313 379 -1307 413
rect -1273 379 -1267 413
rect -1313 341 -1267 379
rect -1313 307 -1307 341
rect -1273 307 -1267 341
rect -1313 269 -1267 307
rect -1313 235 -1307 269
rect -1273 235 -1267 269
rect -1313 197 -1267 235
rect -1313 163 -1307 197
rect -1273 163 -1267 197
rect -1313 125 -1267 163
rect -1313 91 -1307 125
rect -1273 91 -1267 125
rect -1313 53 -1267 91
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -91 -1267 -53
rect -1313 -125 -1307 -91
rect -1273 -125 -1267 -91
rect -1313 -163 -1267 -125
rect -1313 -197 -1307 -163
rect -1273 -197 -1267 -163
rect -1313 -235 -1267 -197
rect -1313 -269 -1307 -235
rect -1273 -269 -1267 -235
rect -1313 -307 -1267 -269
rect -1313 -341 -1307 -307
rect -1273 -341 -1267 -307
rect -1313 -379 -1267 -341
rect -1313 -413 -1307 -379
rect -1273 -413 -1267 -379
rect -1313 -451 -1267 -413
rect -1313 -485 -1307 -451
rect -1273 -485 -1267 -451
rect -1313 -523 -1267 -485
rect -1313 -557 -1307 -523
rect -1273 -557 -1267 -523
rect -1313 -595 -1267 -557
rect -1313 -629 -1307 -595
rect -1273 -629 -1267 -595
rect -1313 -667 -1267 -629
rect -1313 -701 -1307 -667
rect -1273 -701 -1267 -667
rect -1313 -739 -1267 -701
rect -1313 -773 -1307 -739
rect -1273 -773 -1267 -739
rect -1313 -800 -1267 -773
rect -1055 773 -1009 800
rect -1055 739 -1049 773
rect -1015 739 -1009 773
rect -1055 701 -1009 739
rect -1055 667 -1049 701
rect -1015 667 -1009 701
rect -1055 629 -1009 667
rect -1055 595 -1049 629
rect -1015 595 -1009 629
rect -1055 557 -1009 595
rect -1055 523 -1049 557
rect -1015 523 -1009 557
rect -1055 485 -1009 523
rect -1055 451 -1049 485
rect -1015 451 -1009 485
rect -1055 413 -1009 451
rect -1055 379 -1049 413
rect -1015 379 -1009 413
rect -1055 341 -1009 379
rect -1055 307 -1049 341
rect -1015 307 -1009 341
rect -1055 269 -1009 307
rect -1055 235 -1049 269
rect -1015 235 -1009 269
rect -1055 197 -1009 235
rect -1055 163 -1049 197
rect -1015 163 -1009 197
rect -1055 125 -1009 163
rect -1055 91 -1049 125
rect -1015 91 -1009 125
rect -1055 53 -1009 91
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -91 -1009 -53
rect -1055 -125 -1049 -91
rect -1015 -125 -1009 -91
rect -1055 -163 -1009 -125
rect -1055 -197 -1049 -163
rect -1015 -197 -1009 -163
rect -1055 -235 -1009 -197
rect -1055 -269 -1049 -235
rect -1015 -269 -1009 -235
rect -1055 -307 -1009 -269
rect -1055 -341 -1049 -307
rect -1015 -341 -1009 -307
rect -1055 -379 -1009 -341
rect -1055 -413 -1049 -379
rect -1015 -413 -1009 -379
rect -1055 -451 -1009 -413
rect -1055 -485 -1049 -451
rect -1015 -485 -1009 -451
rect -1055 -523 -1009 -485
rect -1055 -557 -1049 -523
rect -1015 -557 -1009 -523
rect -1055 -595 -1009 -557
rect -1055 -629 -1049 -595
rect -1015 -629 -1009 -595
rect -1055 -667 -1009 -629
rect -1055 -701 -1049 -667
rect -1015 -701 -1009 -667
rect -1055 -739 -1009 -701
rect -1055 -773 -1049 -739
rect -1015 -773 -1009 -739
rect -1055 -800 -1009 -773
rect -797 773 -751 800
rect -797 739 -791 773
rect -757 739 -751 773
rect -797 701 -751 739
rect -797 667 -791 701
rect -757 667 -751 701
rect -797 629 -751 667
rect -797 595 -791 629
rect -757 595 -751 629
rect -797 557 -751 595
rect -797 523 -791 557
rect -757 523 -751 557
rect -797 485 -751 523
rect -797 451 -791 485
rect -757 451 -751 485
rect -797 413 -751 451
rect -797 379 -791 413
rect -757 379 -751 413
rect -797 341 -751 379
rect -797 307 -791 341
rect -757 307 -751 341
rect -797 269 -751 307
rect -797 235 -791 269
rect -757 235 -751 269
rect -797 197 -751 235
rect -797 163 -791 197
rect -757 163 -751 197
rect -797 125 -751 163
rect -797 91 -791 125
rect -757 91 -751 125
rect -797 53 -751 91
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -91 -751 -53
rect -797 -125 -791 -91
rect -757 -125 -751 -91
rect -797 -163 -751 -125
rect -797 -197 -791 -163
rect -757 -197 -751 -163
rect -797 -235 -751 -197
rect -797 -269 -791 -235
rect -757 -269 -751 -235
rect -797 -307 -751 -269
rect -797 -341 -791 -307
rect -757 -341 -751 -307
rect -797 -379 -751 -341
rect -797 -413 -791 -379
rect -757 -413 -751 -379
rect -797 -451 -751 -413
rect -797 -485 -791 -451
rect -757 -485 -751 -451
rect -797 -523 -751 -485
rect -797 -557 -791 -523
rect -757 -557 -751 -523
rect -797 -595 -751 -557
rect -797 -629 -791 -595
rect -757 -629 -751 -595
rect -797 -667 -751 -629
rect -797 -701 -791 -667
rect -757 -701 -751 -667
rect -797 -739 -751 -701
rect -797 -773 -791 -739
rect -757 -773 -751 -739
rect -797 -800 -751 -773
rect -539 773 -493 800
rect -539 739 -533 773
rect -499 739 -493 773
rect -539 701 -493 739
rect -539 667 -533 701
rect -499 667 -493 701
rect -539 629 -493 667
rect -539 595 -533 629
rect -499 595 -493 629
rect -539 557 -493 595
rect -539 523 -533 557
rect -499 523 -493 557
rect -539 485 -493 523
rect -539 451 -533 485
rect -499 451 -493 485
rect -539 413 -493 451
rect -539 379 -533 413
rect -499 379 -493 413
rect -539 341 -493 379
rect -539 307 -533 341
rect -499 307 -493 341
rect -539 269 -493 307
rect -539 235 -533 269
rect -499 235 -493 269
rect -539 197 -493 235
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -163 -493 -125
rect -539 -197 -533 -163
rect -499 -197 -493 -163
rect -539 -235 -493 -197
rect -539 -269 -533 -235
rect -499 -269 -493 -235
rect -539 -307 -493 -269
rect -539 -341 -533 -307
rect -499 -341 -493 -307
rect -539 -379 -493 -341
rect -539 -413 -533 -379
rect -499 -413 -493 -379
rect -539 -451 -493 -413
rect -539 -485 -533 -451
rect -499 -485 -493 -451
rect -539 -523 -493 -485
rect -539 -557 -533 -523
rect -499 -557 -493 -523
rect -539 -595 -493 -557
rect -539 -629 -533 -595
rect -499 -629 -493 -595
rect -539 -667 -493 -629
rect -539 -701 -533 -667
rect -499 -701 -493 -667
rect -539 -739 -493 -701
rect -539 -773 -533 -739
rect -499 -773 -493 -739
rect -539 -800 -493 -773
rect -281 773 -235 800
rect -281 739 -275 773
rect -241 739 -235 773
rect -281 701 -235 739
rect -281 667 -275 701
rect -241 667 -235 701
rect -281 629 -235 667
rect -281 595 -275 629
rect -241 595 -235 629
rect -281 557 -235 595
rect -281 523 -275 557
rect -241 523 -235 557
rect -281 485 -235 523
rect -281 451 -275 485
rect -241 451 -235 485
rect -281 413 -235 451
rect -281 379 -275 413
rect -241 379 -235 413
rect -281 341 -235 379
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -451 -235 -413
rect -281 -485 -275 -451
rect -241 -485 -235 -451
rect -281 -523 -235 -485
rect -281 -557 -275 -523
rect -241 -557 -235 -523
rect -281 -595 -235 -557
rect -281 -629 -275 -595
rect -241 -629 -235 -595
rect -281 -667 -235 -629
rect -281 -701 -275 -667
rect -241 -701 -235 -667
rect -281 -739 -235 -701
rect -281 -773 -275 -739
rect -241 -773 -235 -739
rect -281 -800 -235 -773
rect -23 773 23 800
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -800 23 -773
rect 235 773 281 800
rect 235 739 241 773
rect 275 739 281 773
rect 235 701 281 739
rect 235 667 241 701
rect 275 667 281 701
rect 235 629 281 667
rect 235 595 241 629
rect 275 595 281 629
rect 235 557 281 595
rect 235 523 241 557
rect 275 523 281 557
rect 235 485 281 523
rect 235 451 241 485
rect 275 451 281 485
rect 235 413 281 451
rect 235 379 241 413
rect 275 379 281 413
rect 235 341 281 379
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -451 281 -413
rect 235 -485 241 -451
rect 275 -485 281 -451
rect 235 -523 281 -485
rect 235 -557 241 -523
rect 275 -557 281 -523
rect 235 -595 281 -557
rect 235 -629 241 -595
rect 275 -629 281 -595
rect 235 -667 281 -629
rect 235 -701 241 -667
rect 275 -701 281 -667
rect 235 -739 281 -701
rect 235 -773 241 -739
rect 275 -773 281 -739
rect 235 -800 281 -773
rect 493 773 539 800
rect 493 739 499 773
rect 533 739 539 773
rect 493 701 539 739
rect 493 667 499 701
rect 533 667 539 701
rect 493 629 539 667
rect 493 595 499 629
rect 533 595 539 629
rect 493 557 539 595
rect 493 523 499 557
rect 533 523 539 557
rect 493 485 539 523
rect 493 451 499 485
rect 533 451 539 485
rect 493 413 539 451
rect 493 379 499 413
rect 533 379 539 413
rect 493 341 539 379
rect 493 307 499 341
rect 533 307 539 341
rect 493 269 539 307
rect 493 235 499 269
rect 533 235 539 269
rect 493 197 539 235
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -163 539 -125
rect 493 -197 499 -163
rect 533 -197 539 -163
rect 493 -235 539 -197
rect 493 -269 499 -235
rect 533 -269 539 -235
rect 493 -307 539 -269
rect 493 -341 499 -307
rect 533 -341 539 -307
rect 493 -379 539 -341
rect 493 -413 499 -379
rect 533 -413 539 -379
rect 493 -451 539 -413
rect 493 -485 499 -451
rect 533 -485 539 -451
rect 493 -523 539 -485
rect 493 -557 499 -523
rect 533 -557 539 -523
rect 493 -595 539 -557
rect 493 -629 499 -595
rect 533 -629 539 -595
rect 493 -667 539 -629
rect 493 -701 499 -667
rect 533 -701 539 -667
rect 493 -739 539 -701
rect 493 -773 499 -739
rect 533 -773 539 -739
rect 493 -800 539 -773
rect 751 773 797 800
rect 751 739 757 773
rect 791 739 797 773
rect 751 701 797 739
rect 751 667 757 701
rect 791 667 797 701
rect 751 629 797 667
rect 751 595 757 629
rect 791 595 797 629
rect 751 557 797 595
rect 751 523 757 557
rect 791 523 797 557
rect 751 485 797 523
rect 751 451 757 485
rect 791 451 797 485
rect 751 413 797 451
rect 751 379 757 413
rect 791 379 797 413
rect 751 341 797 379
rect 751 307 757 341
rect 791 307 797 341
rect 751 269 797 307
rect 751 235 757 269
rect 791 235 797 269
rect 751 197 797 235
rect 751 163 757 197
rect 791 163 797 197
rect 751 125 797 163
rect 751 91 757 125
rect 791 91 797 125
rect 751 53 797 91
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -91 797 -53
rect 751 -125 757 -91
rect 791 -125 797 -91
rect 751 -163 797 -125
rect 751 -197 757 -163
rect 791 -197 797 -163
rect 751 -235 797 -197
rect 751 -269 757 -235
rect 791 -269 797 -235
rect 751 -307 797 -269
rect 751 -341 757 -307
rect 791 -341 797 -307
rect 751 -379 797 -341
rect 751 -413 757 -379
rect 791 -413 797 -379
rect 751 -451 797 -413
rect 751 -485 757 -451
rect 791 -485 797 -451
rect 751 -523 797 -485
rect 751 -557 757 -523
rect 791 -557 797 -523
rect 751 -595 797 -557
rect 751 -629 757 -595
rect 791 -629 797 -595
rect 751 -667 797 -629
rect 751 -701 757 -667
rect 791 -701 797 -667
rect 751 -739 797 -701
rect 751 -773 757 -739
rect 791 -773 797 -739
rect 751 -800 797 -773
rect 1009 773 1055 800
rect 1009 739 1015 773
rect 1049 739 1055 773
rect 1009 701 1055 739
rect 1009 667 1015 701
rect 1049 667 1055 701
rect 1009 629 1055 667
rect 1009 595 1015 629
rect 1049 595 1055 629
rect 1009 557 1055 595
rect 1009 523 1015 557
rect 1049 523 1055 557
rect 1009 485 1055 523
rect 1009 451 1015 485
rect 1049 451 1055 485
rect 1009 413 1055 451
rect 1009 379 1015 413
rect 1049 379 1055 413
rect 1009 341 1055 379
rect 1009 307 1015 341
rect 1049 307 1055 341
rect 1009 269 1055 307
rect 1009 235 1015 269
rect 1049 235 1055 269
rect 1009 197 1055 235
rect 1009 163 1015 197
rect 1049 163 1055 197
rect 1009 125 1055 163
rect 1009 91 1015 125
rect 1049 91 1055 125
rect 1009 53 1055 91
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -91 1055 -53
rect 1009 -125 1015 -91
rect 1049 -125 1055 -91
rect 1009 -163 1055 -125
rect 1009 -197 1015 -163
rect 1049 -197 1055 -163
rect 1009 -235 1055 -197
rect 1009 -269 1015 -235
rect 1049 -269 1055 -235
rect 1009 -307 1055 -269
rect 1009 -341 1015 -307
rect 1049 -341 1055 -307
rect 1009 -379 1055 -341
rect 1009 -413 1015 -379
rect 1049 -413 1055 -379
rect 1009 -451 1055 -413
rect 1009 -485 1015 -451
rect 1049 -485 1055 -451
rect 1009 -523 1055 -485
rect 1009 -557 1015 -523
rect 1049 -557 1055 -523
rect 1009 -595 1055 -557
rect 1009 -629 1015 -595
rect 1049 -629 1055 -595
rect 1009 -667 1055 -629
rect 1009 -701 1015 -667
rect 1049 -701 1055 -667
rect 1009 -739 1055 -701
rect 1009 -773 1015 -739
rect 1049 -773 1055 -739
rect 1009 -800 1055 -773
rect 1267 773 1313 800
rect 1267 739 1273 773
rect 1307 739 1313 773
rect 1267 701 1313 739
rect 1267 667 1273 701
rect 1307 667 1313 701
rect 1267 629 1313 667
rect 1267 595 1273 629
rect 1307 595 1313 629
rect 1267 557 1313 595
rect 1267 523 1273 557
rect 1307 523 1313 557
rect 1267 485 1313 523
rect 1267 451 1273 485
rect 1307 451 1313 485
rect 1267 413 1313 451
rect 1267 379 1273 413
rect 1307 379 1313 413
rect 1267 341 1313 379
rect 1267 307 1273 341
rect 1307 307 1313 341
rect 1267 269 1313 307
rect 1267 235 1273 269
rect 1307 235 1313 269
rect 1267 197 1313 235
rect 1267 163 1273 197
rect 1307 163 1313 197
rect 1267 125 1313 163
rect 1267 91 1273 125
rect 1307 91 1313 125
rect 1267 53 1313 91
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -91 1313 -53
rect 1267 -125 1273 -91
rect 1307 -125 1313 -91
rect 1267 -163 1313 -125
rect 1267 -197 1273 -163
rect 1307 -197 1313 -163
rect 1267 -235 1313 -197
rect 1267 -269 1273 -235
rect 1307 -269 1313 -235
rect 1267 -307 1313 -269
rect 1267 -341 1273 -307
rect 1307 -341 1313 -307
rect 1267 -379 1313 -341
rect 1267 -413 1273 -379
rect 1307 -413 1313 -379
rect 1267 -451 1313 -413
rect 1267 -485 1273 -451
rect 1307 -485 1313 -451
rect 1267 -523 1313 -485
rect 1267 -557 1273 -523
rect 1307 -557 1313 -523
rect 1267 -595 1313 -557
rect 1267 -629 1273 -595
rect 1307 -629 1313 -595
rect 1267 -667 1313 -629
rect 1267 -701 1273 -667
rect 1307 -701 1313 -667
rect 1267 -739 1313 -701
rect 1267 -773 1273 -739
rect 1307 -773 1313 -739
rect 1267 -800 1313 -773
rect -1257 -847 -1065 -841
rect -1257 -881 -1214 -847
rect -1180 -881 -1142 -847
rect -1108 -881 -1065 -847
rect -1257 -887 -1065 -881
rect -999 -847 -807 -841
rect -999 -881 -956 -847
rect -922 -881 -884 -847
rect -850 -881 -807 -847
rect -999 -887 -807 -881
rect -741 -847 -549 -841
rect -741 -881 -698 -847
rect -664 -881 -626 -847
rect -592 -881 -549 -847
rect -741 -887 -549 -881
rect -483 -847 -291 -841
rect -483 -881 -440 -847
rect -406 -881 -368 -847
rect -334 -881 -291 -847
rect -483 -887 -291 -881
rect -225 -847 -33 -841
rect -225 -881 -182 -847
rect -148 -881 -110 -847
rect -76 -881 -33 -847
rect -225 -887 -33 -881
rect 33 -847 225 -841
rect 33 -881 76 -847
rect 110 -881 148 -847
rect 182 -881 225 -847
rect 33 -887 225 -881
rect 291 -847 483 -841
rect 291 -881 334 -847
rect 368 -881 406 -847
rect 440 -881 483 -847
rect 291 -887 483 -881
rect 549 -847 741 -841
rect 549 -881 592 -847
rect 626 -881 664 -847
rect 698 -881 741 -847
rect 549 -887 741 -881
rect 807 -847 999 -841
rect 807 -881 850 -847
rect 884 -881 922 -847
rect 956 -881 999 -847
rect 807 -887 999 -881
rect 1065 -847 1257 -841
rect 1065 -881 1108 -847
rect 1142 -881 1180 -847
rect 1214 -881 1257 -847
rect 1065 -887 1257 -881
<< properties >>
string FIXED_BBOX -1404 -966 1404 966
<< end >>
