** sch_path: /home/ttuser/tt10-DAC-main/xschem/untitled-3.sch
**.subckt untitled-3 OUT OUT_parax
*.opin OUT
*.opin OUT_parax
Vref net4 GND 1.8
V0 D0 GND PULSE(1.8 0 1n 100p 100p 10u 20u)
V1 D2 GND PULSE(1.8 0 1n 100p 100p 40u 80u)
V3 D3 GND PULSE(1.8 0 1n 100p 100p 80u 160u)
V4 D1 GND PULSE(1.8 0 1n 100p 100p 20u 40u)
Vref1 net2 GND 1.8
x1 D3 D2 D0 D1 net4 net5 net1 net3 DAC
Vmeas net2 net1 0
.save i(vmeas)
Vref2 net3 GND 0
R1 OUT net5 500 m=1
C1 net5 GND 5p m=1
Vref3 net9 GND 1.8
V2 D0 GND PULSE(1.8 0 1n 100p 100p 10u 20u)
V5 D2 GND PULSE(1.8 0 1n 100p 100p 40u 80u)
V6 D3 GND PULSE(1.8 0 1n 100p 100p 80u 160u)
V7 D1 GND PULSE(1.8 0 1n 100p 100p 20u 40u)
Vref4 net7 GND 1.8
x2 D3 D2 D0 D1 net9 net10 net6 net8 DAC_parax
Vmeas1 net7 net6 0
.save i(vmeas1)
Vref5 net8 GND 0
R2 OUT_parax net10 500 m=1
C2 net10 GND 5p m=1
**** begin user architecture code



.option savecurrents
.control
save all
  op
  remzerovec
  write untitled-3.raw
  set appendwrite
  tran 2n 160u
  remzerovec
  write untitled-3.raw
  set appendwrite

.endc




** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  DAC.sym # of pins=8
** sym_path: /home/ttuser/tt10-DAC-main/xschem/DAC.sym
** sch_path: /home/ttuser/tt10-DAC-main/xschem/DAC.sch
.subckt DAC D3 D2 D0 D1 Vref OUT VDD VSS
*.ipin D0
*.ipin D1
*.ipin D2
*.ipin D3
*.iopin Vref
*.opin OUT
*.iopin VDD
*.iopin VSS
XR3 net5 Vref VSS sky130_fd_pr__res_xhigh_po_0p35 L=16 mult=1 m=1
XR4 G net5 VSS sky130_fd_pr__res_xhigh_po_0p35 L=16 mult=1 m=1
XR5 VDD OUT VSS sky130_fd_pr__res_xhigh_po_0p69 L=1.75 mult=1 m=1
XM6 OUT D0 net4 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=6 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 OUT D1 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=6 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT D2 net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=6 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT D3 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=6 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 G G VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=8 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 G VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=8 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 G VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=16 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 G VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=33 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net3 G VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.18 W=69 nf=24 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  DAC_parax.sym # of pins=8
** sym_path: /home/ttuser/tt10-DAC-main/xschem/DAC.sym
* NGSPICE file created from DAC_parax.ext - technology: sky130A

.subckt DAC_parax D3 D2 D0 D1 Vref OUT VDD VSS
X0 a_3992_n1502# D2.t0 OUT.t12 VSS.t107 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.59 ps=4.59 w=2 l=0.18
X1 OUT.t11 D2.t1 a_3992_n1502# VSS.t106 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.18
X2 a_3992_n1502# D2.t2 OUT.t10 VSS.t105 sky130_fd_pr__nfet_01v8_lvt ad=0.59 pd=4.59 as=0.3 ps=2.3 w=2 l=0.18
X3 VSS.t71 a_n1186_n1046.t7 a_1632_n1418# VSS.t70 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.78765 ps=5.93 w=2.67 l=0.18
X4 VSS.t36 a_n1186_n1046.t8 a_2756_n1382# VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X5 VSS.t85 a_n1186_n1046.t9 a_5585_876.t26 VSS.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X6 a_n1774_2554# a_n1186_n1046.t6 VSS.t108 sky130_fd_pr__res_xhigh_po_0p35 l=16
X7 VSS.t73 a_n1186_n1046.t4 a_n1186_n1046.t5 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.78765 ps=5.93 w=2.67 l=0.18
X8 a_5585_876.t25 a_n1186_n1046.t10 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X9 VSS.t34 a_n1186_n1046.t11 a_5585_876.t24 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X10 a_2756_n1382# a_n1186_n1046.t12 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X11 VSS.t7 a_n1186_n1046.t13 a_2756_n1382# VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X12 a_5585_876.t23 a_n1186_n1046.t14 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X13 a_5585_876.t22 a_n1186_n1046.t15 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X14 a_n1186_n1046.t3 a_n1186_n1046.t2 VSS.t87 VSS.t86 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X15 VSS.t83 a_n1186_n1046.t16 a_5585_876.t21 VSS.t82 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X16 a_5585_876.t20 a_n1186_n1046.t17 VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X17 a_5585_876.t19 a_n1186_n1046.t18 VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X18 a_3992_n1502# a_n1186_n1046.t19 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X19 VSS.t102 a_n1186_n1046.t20 a_5585_876.t18 VSS.t101 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X20 a_1632_n1418# D0.t0 OUT.t6 VSS.t90 sky130_fd_pr__nfet_01v8_lvt ad=0.59 pd=4.59 as=0.3 ps=2.3 w=2 l=0.18
X21 a_2756_n1382# a_n1186_n1046.t21 VSS.t96 VSS.t95 sky130_fd_pr__nfet_01v8_lvt ad=0.78765 pd=5.93 as=0.4005 ps=2.97 w=2.67 l=0.18
X22 VSS.t26 a_n1186_n1046.t22 a_3992_n1502# VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X23 a_1632_n1418# D0.t1 OUT.t5 VSS.t89 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.59 ps=4.59 w=2 l=0.18
X24 OUT.t4 D0.t2 a_1632_n1418# VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.18
X25 VSS.t100 a_n1186_n1046.t23 a_5585_876.t17 VSS.t99 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X26 VSS.t94 a_n1186_n1046.t24 a_5585_876.t16 VSS.t93 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X27 VSS.t10 a_n1186_n1046.t25 a_3992_n1502# VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X28 a_5585_876.t15 a_n1186_n1046.t26 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X29 a_5585_876.t2 D3.t0 OUT.t9 VSS.t104 sky130_fd_pr__nfet_01v8_lvt ad=0.59 pd=4.59 as=0.3 ps=2.3 w=2 l=0.18
X30 a_1632_n1418# a_n1186_n1046.t27 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X31 a_3992_n1502# a_n1186_n1046.t28 VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X32 VSS.t42 a_n1186_n1046.t29 a_3992_n1502# VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X33 a_n1774_2554# Vref.t0 VSS.t92 sky130_fd_pr__res_xhigh_po_0p35 l=16
X34 a_5585_876.t1 D3.t1 OUT.t8 VSS.t103 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.59 ps=4.59 w=2 l=0.18
X35 OUT.t3 D3.t2 a_5585_876.t0 VSS.t81 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.18
X36 a_5585_876.t14 a_n1186_n1046.t30 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X37 VSS.t16 a_n1186_n1046.t31 a_3992_n1502# VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.81125 ps=6.09 w=2.75 l=0.18
X38 a_3992_n1502# a_n1186_n1046.t32 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X39 VSS.t61 a_n1186_n1046.t33 a_1632_n1418# VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=0.78765 pd=5.93 as=0.4005 ps=2.97 w=2.67 l=0.18
X40 VSS.t30 a_n1186_n1046.t34 a_5585_876.t13 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X41 VSS.t65 a_n1186_n1046.t0 a_n1186_n1046.t1 VSS.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.78765 pd=5.93 as=0.4005 ps=2.97 w=2.67 l=0.18
X42 OUT.t7 VDD.t0 VSS.t91 sky130_fd_pr__res_xhigh_po_0p69 l=1.75
X43 OUT.t0 D1.t0 a_2756_n1382# VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.18
X44 a_2756_n1382# D1.t1 OUT.t1 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.59 pd=4.59 as=0.3 ps=2.3 w=2 l=0.18
X45 a_5585_876.t12 a_n1186_n1046.t35 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X46 VSS.t80 a_n1186_n1046.t36 a_2756_n1382# VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.78765 ps=5.93 w=2.67 l=0.18
X47 VSS.t38 a_n1186_n1046.t37 a_5585_876.t11 VSS.t37 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.8496 ps=6.35 w=2.88 l=0.18
X48 a_5585_876.t10 a_n1186_n1046.t38 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X49 VSS.t59 a_n1186_n1046.t39 a_5585_876.t9 VSS.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X50 VSS.t110 a_n1186_n1046.t40 a_5585_876.t8 VSS.t109 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X51 a_5585_876.t7 a_n1186_n1046.t41 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.8496 pd=6.35 as=0.432 ps=3.18 w=2.88 l=0.18
X52 a_3992_n1502# a_n1186_n1046.t42 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.81125 pd=6.09 as=0.4125 ps=3.05 w=2.75 l=0.18
X53 VSS.t5 a_n1186_n1046.t43 a_5585_876.t6 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X54 a_5585_876.t5 a_n1186_n1046.t44 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X55 a_2756_n1382# a_n1186_n1046.t45 VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X56 a_3992_n1502# a_n1186_n1046.t46 VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X57 a_5585_876.t4 a_n1186_n1046.t47 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X58 VSS.t78 a_n1186_n1046.t48 a_5585_876.t3 VSS.t77 sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X59 VSS.t98 a_n1186_n1046.t49 a_3992_n1502# VSS.t97 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X60 a_2756_n1382# D1.t2 OUT.t2 VSS.t74 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.59 ps=4.59 w=2 l=0.18
X61 VSS.t57 a_n1186_n1046.t50 a_3992_n1502# VSS.t56 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X62 a_3992_n1502# a_n1186_n1046.t51 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
R0 D2.n1 D2.t1 483.647
R1 D2.n0 D2.t0 483.113
R2 D2.n0 D2.t2 482.634
R3 D2 D2.n1 5.65562
R4 D2.n1 D2.n0 1.99752
R5 OUT.n3 OUT.n2 42.6841
R6 OUT.n1 OUT.n0 42.659
R7 OUT.n9 OUT.n8 42.6109
R8 OUT.n5 OUT.n4 42.4848
R9 OUT.n9 OUT.t8 42.0916
R10 OUT.n1 OUT.t12 42.0807
R11 OUT.n3 OUT.t2 41.9969
R12 OUT.n5 OUT.t5 41.9058
R13 OUT.n11 OUT.t7 22.8927
R14 OUT.n4 OUT.t6 9.0005
R15 OUT.n4 OUT.t4 9.0005
R16 OUT.n2 OUT.t1 9.0005
R17 OUT.n2 OUT.t0 9.0005
R18 OUT.n0 OUT.t10 9.0005
R19 OUT.n0 OUT.t11 9.0005
R20 OUT.n8 OUT.t9 9.0005
R21 OUT.n8 OUT.t3 9.0005
R22 OUT.n6 OUT.n5 5.65959
R23 OUT.n7 OUT.n6 3.75902
R24 OUT.n10 OUT.n7 3.59425
R25 OUT.n11 OUT.n10 3.38402
R26 OUT.n6 OUT.n3 2.17312
R27 OUT.n7 OUT.n1 2.14633
R28 OUT.n10 OUT.n9 1.9217
R29 OUT OUT.n11 0.207578
R30 VSS.n34 VSS.n26 13094.7
R31 VSS.n29 VSS.n26 13094.7
R32 VSS.n34 VSS.n27 13094.7
R33 VSS.n38 VSS.n21 13094.7
R34 VSS.n38 VSS.n22 13094.7
R35 VSS.n39 VSS.n21 13094.7
R36 VSS.n39 VSS.n22 13094.7
R37 VSS.n136 VSS.n96 9815.24
R38 VSS.n136 VSS.n97 9815.24
R39 VSS.n138 VSS.n96 9815.24
R40 VSS.n138 VSS.n97 9815.24
R41 VSS.n121 VSS.n67 6402.5
R42 VSS.n158 VSS.n67 6402.5
R43 VSS.n121 VSS.n68 6402.5
R44 VSS.n158 VSS.n68 6402.5
R45 VSS.n102 VSS.n98 5035.09
R46 VSS.n133 VSS.n98 5035.09
R47 VSS.n102 VSS.n99 5035.09
R48 VSS.n133 VSS.n99 5035.09
R49 VSS.n164 VSS.n64 4687.44
R50 VSS.n169 VSS.n64 4687.44
R51 VSS.n164 VSS.n65 4687.44
R52 VSS.n169 VSS.n65 4687.44
R53 VSS.n182 VSS.n14 3853.09
R54 VSS.n23 VSS.n14 3853.09
R55 VSS.n182 VSS.n15 3853.09
R56 VSS.n23 VSS.n15 3853.09
R57 VSS.n53 VSS.n11 3853.09
R58 VSS.n185 VSS.n11 3853.09
R59 VSS.n53 VSS.n12 3853.09
R60 VSS.n185 VSS.n12 3853.09
R61 VSS.n125 VSS.n106 3464.88
R62 VSS.n125 VSS.n107 3464.88
R63 VSS.n126 VSS.n106 3464.88
R64 VSS.n126 VSS.n107 3464.88
R65 VSS.n62 VSS.n55 3464.88
R66 VSS.n57 VSS.n55 3464.88
R67 VSS.n62 VSS.n56 3464.88
R68 VSS.n57 VSS.n56 3464.88
R69 VSS.n161 VSS.n51 3464.88
R70 VSS.n172 VSS.n51 3464.88
R71 VSS.n161 VSS.n49 3464.88
R72 VSS.n172 VSS.n49 3464.88
R73 VSS.n119 VSS.n111 3464.88
R74 VSS.n115 VSS.n111 3464.88
R75 VSS.n119 VSS.n112 3464.88
R76 VSS.n115 VSS.n112 3464.88
R77 VSS.n37 VSS.n20 850.823
R78 VSS.n37 VSS.n19 850.823
R79 VSS.n31 VSS.n30 850.823
R80 VSS.n33 VSS.n31 850.823
R81 VSS.n40 VSS.n20 838.206
R82 VSS.n33 VSS.n32 837.894
R83 VSS.n30 VSS.n18 837.361
R84 VSS.n41 VSS.n19 836.61
R85 VSS.n25 VSS.n24 825.288
R86 VSS.n184 VSS.n183 737.688
R87 VSS.n135 VSS.n95 637.741
R88 VSS.n135 VSS.n94 637.741
R89 VSS.n170 VSS.n63 453.372
R90 VSS.n70 VSS.n69 416
R91 VSS.n157 VSS.n69 416
R92 VSS.n139 VSS.n95 405.986
R93 VSS.n140 VSS.n94 404.276
R94 VSS.n157 VSS.n156 335.334
R95 VSS.n155 VSS.n70 334.32
R96 VSS.n163 VSS.n159 331.959
R97 VSS.n132 VSS.n100 327.154
R98 VSS.n103 VSS.n100 327.154
R99 VSS.n165 VSS.n66 304.565
R100 VSS.n168 VSS.n66 304.565
R101 VSS.n40 VSS.n39 292.5
R102 VSS.n39 VSS.t108 292.5
R103 VSS.n38 VSS.n37 292.5
R104 VSS.t108 VSS.n38 292.5
R105 VSS.n32 VSS.n27 292.5
R106 VSS.n31 VSS.n26 292.5
R107 VSS.n26 VSS.t92 292.5
R108 VSS.n28 VSS.n27 283.495
R109 VSS.n168 VSS.n167 261.43
R110 VSS.n166 VSS.n165 258.897
R111 VSS.n181 VSS.n16 250.353
R112 VSS.n17 VSS.n16 250.353
R113 VSS.n52 VSS.n10 250.353
R114 VSS.n186 VSS.n10 250.353
R115 VSS.n52 VSS.n9 226.244
R116 VSS.n187 VSS.n186 225.232
R117 VSS.n173 VSS.n50 225.13
R118 VSS.n50 VSS.n48 225.13
R119 VSS.n116 VSS.n113 225.13
R120 VSS.n118 VSS.n113 225.13
R121 VSS.n124 VSS.n105 225.13
R122 VSS.n124 VSS.n104 225.13
R123 VSS.n59 VSS.n58 225.13
R124 VSS.n61 VSS.n59 225.13
R125 VSS.n36 VSS.n35 224.381
R126 VSS.n181 VSS.n180 221.222
R127 VSS.n179 VSS.n17 220.157
R128 VSS.n132 VSS.n131 215.095
R129 VSS.n130 VSS.n103 212.882
R130 VSS.n127 VSS.n105 206.962
R131 VSS.n174 VSS.n173 206.371
R132 VSS.n117 VSS.n116 206.371
R133 VSS.n174 VSS.n48 206.371
R134 VSS.n118 VSS.n117 206.371
R135 VSS.n128 VSS.n104 204.113
R136 VSS.n61 VSS.n60 202.843
R137 VSS.n58 VSS.n46 201.352
R138 VSS.n102 VSS.n101 199.612
R139 VSS.n133 VSS.n132 195
R140 VSS.n134 VSS.n133 195
R141 VSS.n103 VSS.n102 195
R142 VSS.n101 VSS.t27 124.486
R143 VSS.t103 VSS.n123 124.486
R144 VSS.n122 VSS.t17 124.486
R145 VSS.n159 VSS.t15 124.486
R146 VSS.n163 VSS.t95 124.486
R147 VSS.n183 VSS.t64 124.486
R148 VSS.n24 VSS.t72 124.486
R149 VSS.n29 VSS.n28 119.677
R150 VSS.n12 VSS.n9 117.001
R151 VSS.t19 VSS.n12 117.001
R152 VSS.n11 VSS.n10 117.001
R153 VSS.t19 VSS.n11 117.001
R154 VSS.n180 VSS.n15 117.001
R155 VSS.t86 VSS.n15 117.001
R156 VSS.n16 VSS.n14 117.001
R157 VSS.t86 VSS.n14 117.001
R158 VSS.n117 VSS.n112 117.001
R159 VSS.t106 VSS.n112 117.001
R160 VSS.n113 VSS.n111 117.001
R161 VSS.t106 VSS.n111 117.001
R162 VSS.n174 VSS.n49 117.001
R163 VSS.t8 VSS.n49 117.001
R164 VSS.n51 VSS.n50 117.001
R165 VSS.t8 VSS.n51 117.001
R166 VSS.n60 VSS.n56 117.001
R167 VSS.n56 VSS.t88 117.001
R168 VSS.n59 VSS.n55 117.001
R169 VSS.t88 VSS.n55 117.001
R170 VSS.n127 VSS.n126 117.001
R171 VSS.n126 VSS.t81 117.001
R172 VSS.n125 VSS.n124 117.001
R173 VSS.t81 VSS.n125 117.001
R174 VSS.t108 VSS.n25 113.728
R175 VSS.t108 VSS.n36 113.728
R176 VSS.n35 VSS.t92 113.728
R177 VSS.t90 VSS.n54 110.653
R178 VSS.t70 VSS.n13 110.653
R179 VSS.n123 VSS.n122 90.6746
R180 VSS.t27 VSS.t109 73.7693
R181 VSS.t109 VSS.t23 73.7693
R182 VSS.t23 VSS.t101 73.7693
R183 VSS.t101 VSS.t0 73.7693
R184 VSS.t0 VSS.t77 73.7693
R185 VSS.t62 VSS.t93 73.7693
R186 VSS.t93 VSS.t68 73.7693
R187 VSS.t68 VSS.t33 73.7693
R188 VSS.t33 VSS.t13 73.7693
R189 VSS.t13 VSS.t4 73.7693
R190 VSS.t43 VSS.t99 73.7693
R191 VSS.t82 VSS.t43 73.7693
R192 VSS.t47 VSS.t82 73.7693
R193 VSS.t58 VSS.t47 73.7693
R194 VSS.t51 VSS.t58 73.7693
R195 VSS.t29 VSS.t51 73.7693
R196 VSS.t45 VSS.t29 73.7693
R197 VSS.t84 VSS.t45 73.7693
R198 VSS.t54 VSS.t84 73.7693
R199 VSS.t81 VSS.t103 73.7693
R200 VSS.t17 VSS.t41 73.7693
R201 VSS.t41 VSS.t21 73.7693
R202 VSS.t21 VSS.t25 73.7693
R203 VSS.t25 VSS.t11 73.7693
R204 VSS.t11 VSS.t97 73.7693
R205 VSS.t9 VSS.t39 73.7693
R206 VSS.t6 VSS.t2 73.7693
R207 VSS.t86 VSS.t64 73.7693
R208 VSS.t72 VSS.t86 73.7693
R209 VSS.n116 VSS.n115 73.1255
R210 VSS.n115 VSS.n114 73.1255
R211 VSS.n119 VSS.n118 73.1255
R212 VSS.n120 VSS.n119 73.1255
R213 VSS.n173 VSS.n172 73.1255
R214 VSS.n172 VSS.n171 73.1255
R215 VSS.n161 VSS.n48 73.1255
R216 VSS.n162 VSS.n161 73.1255
R217 VSS.n58 VSS.n57 73.1255
R218 VSS.n57 VSS.n13 73.1255
R219 VSS.n62 VSS.n61 73.1255
R220 VSS.n63 VSS.n62 73.1255
R221 VSS.n107 VSS.n105 73.1255
R222 VSS.n123 VSS.n107 73.1255
R223 VSS.n106 VSS.n104 73.1255
R224 VSS.n108 VSS.n106 73.1255
R225 VSS.t104 VSS.t37 72.2324
R226 VSS.t66 VSS.t105 72.2324
R227 VSS.t56 VSS.t106 72.2324
R228 VSS.t75 VSS.t107 72.2324
R229 VSS.t8 VSS.t49 72.2324
R230 VSS.t74 VSS.t79 72.2324
R231 VSS.n171 VSS.n170 72.2324
R232 VSS.t31 VSS.n134 67.6219
R233 VSS.t88 VSS.t60 59.9376
R234 VSS.t19 VSS.t89 59.9376
R235 VSS.n158 VSS.n157 58.5005
R236 VSS.n159 VSS.n158 58.5005
R237 VSS.n121 VSS.n70 58.5005
R238 VSS.n122 VSS.n121 58.5005
R239 VSS.n186 VSS.n185 58.5005
R240 VSS.n185 VSS.n184 58.5005
R241 VSS.n53 VSS.n52 58.5005
R242 VSS.n54 VSS.n53 58.5005
R243 VSS.n169 VSS.n168 58.5005
R244 VSS.n170 VSS.n169 58.5005
R245 VSS.n167 VSS.n65 58.5005
R246 VSS.n160 VSS.n65 58.5005
R247 VSS.n165 VSS.n164 58.5005
R248 VSS.n164 VSS.n163 58.5005
R249 VSS.n66 VSS.n64 58.5005
R250 VSS.n160 VSS.n64 58.5005
R251 VSS.n23 VSS.n17 58.5005
R252 VSS.n24 VSS.n23 58.5005
R253 VSS.n182 VSS.n181 58.5005
R254 VSS.n183 VSS.n182 58.5005
R255 VSS.n97 VSS.n95 53.1823
R256 VSS.n109 VSS.n97 53.1823
R257 VSS.n96 VSS.n94 53.1823
R258 VSS.n101 VSS.n96 53.1823
R259 VSS.t37 VSS.n108 52.2534
R260 VSS.n109 VSS.t104 52.2534
R261 VSS.n114 VSS.t75 52.2534
R262 VSS.n171 VSS.t79 52.2534
R263 VSS.n162 VSS.t6 49.1797
R264 VSS.t77 VSS.t91 43.0323
R265 VSS.n137 VSS.t4 36.8849
R266 VSS.n137 VSS.t31 36.8849
R267 VSS.t39 VSS.n110 36.8849
R268 VSS.n160 VSS.t35 36.8849
R269 VSS.n44 VSS.t65 36.7226
R270 VSS.n7 VSS.t61 36.7169
R271 VSS.t53 VSS.n160 35.348
R272 VSS.n156 VSS.n68 32.5005
R273 VSS.n110 VSS.n68 32.5005
R274 VSS.n69 VSS.n67 32.5005
R275 VSS.n110 VSS.n67 32.5005
R276 VSS.n131 VSS.n99 32.5005
R277 VSS.t91 VSS.n99 32.5005
R278 VSS.n100 VSS.n98 32.5005
R279 VSS.t91 VSS.n98 32.5005
R280 VSS.t91 VSS.t62 30.7375
R281 VSS.n3 VSS.n1 29.9991
R282 VSS.n73 VSS.n71 29.9799
R283 VSS.n144 VSS.n142 29.9715
R284 VSS.n152 VSS.n151 29.5696
R285 VSS.n150 VSS.n149 29.5588
R286 VSS.n148 VSS.n147 29.5479
R287 VSS.n146 VSS.n145 29.5425
R288 VSS.n144 VSS.n143 29.537
R289 VSS.n5 VSS.n4 29.5207
R290 VSS.n7 VSS.n6 29.5153
R291 VSS.n3 VSS.n2 29.5153
R292 VSS.n44 VSS.n43 29.5098
R293 VSS.n73 VSS.n72 29.4498
R294 VSS.n89 VSS.n88 29.4443
R295 VSS.n75 VSS.n74 29.4443
R296 VSS.n81 VSS.n80 29.4389
R297 VSS.n77 VSS.n76 29.4389
R298 VSS.n87 VSS.n86 29.4334
R299 VSS.n83 VSS.n82 29.4334
R300 VSS.n79 VSS.n78 29.4334
R301 VSS.n93 VSS.n92 29.428
R302 VSS.n91 VSS.n90 29.428
R303 VSS.n85 VSS.n84 29.428
R304 VSS.t97 VSS.n120 24.5901
R305 VSS.t95 VSS.n162 24.5901
R306 VSS.n108 VSS.t54 21.5164
R307 VSS.t81 VSS.n109 21.5164
R308 VSS.n114 VSS.t15 21.5164
R309 VSS.n136 VSS.n135 16.7148
R310 VSS.n137 VSS.n136 16.7148
R311 VSS.n139 VSS.n138 16.7148
R312 VSS.n138 VSS.n137 16.7148
R313 VSS.n63 VSS.n54 13.8321
R314 VSS.t60 VSS.t90 13.8321
R315 VSS.t88 VSS.t19 13.8321
R316 VSS.t89 VSS.t70 13.8321
R317 VSS.n184 VSS.n13 13.8321
R318 VSS.n120 VSS.n110 12.2953
R319 VSS.n177 VSS.n176 10.1753
R320 VSS.n22 VSS.n20 9.7505
R321 VSS.n36 VSS.n22 9.7505
R322 VSS.n21 VSS.n19 9.7505
R323 VSS.n25 VSS.n21 9.7505
R324 VSS.n30 VSS.n29 9.7505
R325 VSS.n34 VSS.n33 9.7505
R326 VSS.n35 VSS.n34 9.7505
R327 VSS.n6 VSS.t20 6.74207
R328 VSS.n6 VSS.t71 6.74207
R329 VSS.n43 VSS.t87 6.74207
R330 VSS.n43 VSS.t73 6.74207
R331 VSS.n4 VSS.t50 6.74207
R332 VSS.n4 VSS.t80 6.74207
R333 VSS.n2 VSS.t3 6.74207
R334 VSS.n2 VSS.t36 6.74207
R335 VSS.n1 VSS.t96 6.74207
R336 VSS.n1 VSS.t7 6.74207
R337 VSS.n129 VSS.n47 6.63797
R338 VSS.n151 VSS.t76 6.54595
R339 VSS.n151 VSS.t16 6.54595
R340 VSS.n149 VSS.t67 6.54595
R341 VSS.n149 VSS.t57 6.54595
R342 VSS.n147 VSS.t40 6.54595
R343 VSS.n147 VSS.t10 6.54595
R344 VSS.n145 VSS.t12 6.54595
R345 VSS.n145 VSS.t98 6.54595
R346 VSS.n143 VSS.t22 6.54595
R347 VSS.n143 VSS.t26 6.54595
R348 VSS.n142 VSS.t18 6.54595
R349 VSS.n142 VSS.t42 6.54595
R350 VSS.n189 VSS.n5 6.51952
R351 VSS.n176 VSS.n46 6.42018
R352 VSS.n175 VSS.n174 6.41272
R353 VSS.n117 VSS.n47 6.38527
R354 VSS.n8 VSS.n7 6.31358
R355 VSS.n92 VSS.t55 6.2505
R356 VSS.n92 VSS.t38 6.2505
R357 VSS.n90 VSS.t46 6.2505
R358 VSS.n90 VSS.t85 6.2505
R359 VSS.n88 VSS.t52 6.2505
R360 VSS.n88 VSS.t30 6.2505
R361 VSS.n86 VSS.t48 6.2505
R362 VSS.n86 VSS.t59 6.2505
R363 VSS.n84 VSS.t44 6.2505
R364 VSS.n84 VSS.t83 6.2505
R365 VSS.n82 VSS.t32 6.2505
R366 VSS.n82 VSS.t100 6.2505
R367 VSS.n80 VSS.t14 6.2505
R368 VSS.n80 VSS.t5 6.2505
R369 VSS.n78 VSS.t69 6.2505
R370 VSS.n78 VSS.t34 6.2505
R371 VSS.n76 VSS.t63 6.2505
R372 VSS.n76 VSS.t94 6.2505
R373 VSS.n74 VSS.t1 6.2505
R374 VSS.n74 VSS.t78 6.2505
R375 VSS.n72 VSS.t24 6.2505
R376 VSS.n72 VSS.t102 6.2505
R377 VSS.n71 VSS.t28 6.2505
R378 VSS.n71 VSS.t110 6.2505
R379 VSS.n134 VSS.t99 6.1479
R380 VSS.n141 VSS.n93 6.06064
R381 VSS.n153 VSS.n152 6.00166
R382 VSS.n45 VSS.n44 5.42623
R383 VSS.n42 VSS.n18 5.21865
R384 VSS.n42 VSS.n41 4.6505
R385 VSS.n130 VSS.n129 4.11587
R386 VSS.n28 VSS.t92 2.67422
R387 VSS.n175 VSS.n47 2.14119
R388 VSS.n179 VSS.n178 2.02066
R389 VSS.n188 VSS.n187 2.01089
R390 VSS.n176 VSS.n175 2.0005
R391 VSS.n129 VSS.n128 1.8605
R392 VSS.n128 VSS.n127 1.67007
R393 VSS.n178 VSS.n45 1.637
R394 VSS.t105 VSS.t9 1.53735
R395 VSS.t106 VSS.t66 1.53735
R396 VSS.t107 VSS.t56 1.53735
R397 VSS.t2 VSS.t53 1.53735
R398 VSS.t35 VSS.t8 1.53735
R399 VSS.t49 VSS.t74 1.53735
R400 VSS.n167 VSS.n166 1.23127
R401 VSS.n166 VSS.n0 1.03383
R402 VSS.n141 VSS.n140 0.892169
R403 VSS.n131 VSS.n130 0.8005
R404 VSS.n60 VSS.n46 0.7685
R405 VSS.n41 VSS.n40 0.662569
R406 VSS.n45 VSS.n42 0.579283
R407 VSS.n140 VSS.n139 0.549071
R408 VSS.n155 VSS.n154 0.547559
R409 VSS.n85 VSS.n83 0.542641
R410 VSS.n75 VSS.n73 0.536062
R411 VSS.n77 VSS.n75 0.536062
R412 VSS.n81 VSS.n79 0.536062
R413 VSS.n83 VSS.n81 0.536062
R414 VSS.n87 VSS.n85 0.536062
R415 VSS.n89 VSS.n87 0.536062
R416 VSS.n91 VSS.n89 0.536062
R417 VSS.n93 VSS.n91 0.536062
R418 VSS.n79 VSS.n77 0.529483
R419 VSS.n5 VSS.n3 0.494708
R420 VSS.n187 VSS.n9 0.492808
R421 VSS.n156 VSS.n155 0.492808
R422 VSS.n148 VSS.n146 0.45081
R423 VSS.n152 VSS.n150 0.45081
R424 VSS.n146 VSS.n144 0.445601
R425 VSS.n180 VSS.n179 0.441879
R426 VSS.n150 VSS.n148 0.440393
R427 VSS.n154 VSS.n141 0.339145
R428 VSS.n154 VSS.n153 0.267471
R429 VSS VSS.n190 0.259272
R430 VSS.n153 VSS.n0 0.25085
R431 VSS.n177 VSS.n8 0.245181
R432 VSS.n189 VSS.n188 0.231883
R433 VSS.n32 VSS.n18 0.22119
R434 VSS.n178 VSS.n177 0.162734
R435 VSS.n190 VSS.n189 0.160961
R436 VSS.n188 VSS.n8 0.113975
R437 VSS.n190 VSS.n0 0.0589449
R438 a_n1186_n1046.n11 a_n1186_n1046.t47 600.937
R439 a_n1186_n1046.n0 a_n1186_n1046.t37 600.883
R440 a_n1186_n1046.n11 a_n1186_n1046.t14 600.457
R441 a_n1186_n1046.n12 a_n1186_n1046.t35 600.457
R442 a_n1186_n1046.n13 a_n1186_n1046.t10 600.457
R443 a_n1186_n1046.n14 a_n1186_n1046.t17 600.457
R444 a_n1186_n1046.n15 a_n1186_n1046.t30 600.457
R445 a_n1186_n1046.n16 a_n1186_n1046.t44 600.457
R446 a_n1186_n1046.n17 a_n1186_n1046.t18 600.457
R447 a_n1186_n1046.n18 a_n1186_n1046.t38 600.457
R448 a_n1186_n1046.n19 a_n1186_n1046.t15 600.457
R449 a_n1186_n1046.n20 a_n1186_n1046.t26 600.457
R450 a_n1186_n1046.n21 a_n1186_n1046.t41 600.457
R451 a_n1186_n1046.n10 a_n1186_n1046.t40 600.457
R452 a_n1186_n1046.n9 a_n1186_n1046.t20 600.457
R453 a_n1186_n1046.n8 a_n1186_n1046.t48 600.457
R454 a_n1186_n1046.n7 a_n1186_n1046.t24 600.457
R455 a_n1186_n1046.n6 a_n1186_n1046.t11 600.457
R456 a_n1186_n1046.n5 a_n1186_n1046.t43 600.457
R457 a_n1186_n1046.n4 a_n1186_n1046.t23 600.457
R458 a_n1186_n1046.n3 a_n1186_n1046.t16 600.457
R459 a_n1186_n1046.n2 a_n1186_n1046.t39 600.457
R460 a_n1186_n1046.n1 a_n1186_n1046.t34 600.457
R461 a_n1186_n1046.n0 a_n1186_n1046.t9 600.457
R462 a_n1186_n1046.n28 a_n1186_n1046.t46 583.577
R463 a_n1186_n1046.n23 a_n1186_n1046.t31 583.553
R464 a_n1186_n1046.n32 a_n1186_n1046.t42 583.051
R465 a_n1186_n1046.n31 a_n1186_n1046.t28 583.051
R466 a_n1186_n1046.n30 a_n1186_n1046.t51 583.051
R467 a_n1186_n1046.n29 a_n1186_n1046.t32 583.051
R468 a_n1186_n1046.n28 a_n1186_n1046.t19 583.051
R469 a_n1186_n1046.n27 a_n1186_n1046.t29 583.051
R470 a_n1186_n1046.n26 a_n1186_n1046.t22 583.051
R471 a_n1186_n1046.n25 a_n1186_n1046.t49 583.051
R472 a_n1186_n1046.n24 a_n1186_n1046.t25 583.051
R473 a_n1186_n1046.n23 a_n1186_n1046.t50 583.051
R474 a_n1186_n1046.n45 a_n1186_n1046.t2 573.937
R475 a_n1186_n1046.n42 a_n1186_n1046.t27 573.548
R476 a_n1186_n1046.n44 a_n1186_n1046.t4 573.096
R477 a_n1186_n1046.n37 a_n1186_n1046.t45 573.056
R478 a_n1186_n1046.n35 a_n1186_n1046.t36 573.024
R479 a_n1186_n1046.n41 a_n1186_n1046.t7 572.875
R480 a_n1186_n1046.n41 a_n1186_n1046.t33 572.34
R481 a_n1186_n1046.n36 a_n1186_n1046.t13 572.34
R482 a_n1186_n1046.n35 a_n1186_n1046.t8 572.34
R483 a_n1186_n1046.n38 a_n1186_n1046.t21 572.34
R484 a_n1186_n1046.n37 a_n1186_n1046.t12 572.34
R485 a_n1186_n1046.n44 a_n1186_n1046.t0 572.34
R486 a_n1186_n1046.n48 a_n1186_n1046.n47 34.5589
R487 a_n1186_n1046.n48 a_n1186_n1046.t5 31.784
R488 a_n1186_n1046.n34 a_n1186_n1046.n22 9.14921
R489 a_n1186_n1046.n47 a_n1186_n1046.t1 6.74207
R490 a_n1186_n1046.n47 a_n1186_n1046.t3 6.74207
R491 a_n1186_n1046.t6 a_n1186_n1046.n49 6.23175
R492 a_n1186_n1046.n40 a_n1186_n1046.n39 5.987
R493 a_n1186_n1046.n34 a_n1186_n1046.n33 5.81806
R494 a_n1186_n1046.n43 a_n1186_n1046.n42 5.67034
R495 a_n1186_n1046.n39 a_n1186_n1046.n36 4.09326
R496 a_n1186_n1046.n45 a_n1186_n1046.n44 4.05252
R497 a_n1186_n1046.n46 a_n1186_n1046.n43 2.95139
R498 a_n1186_n1046.n49 a_n1186_n1046.n46 2.8855
R499 a_n1186_n1046.n33 a_n1186_n1046.n27 2.80523
R500 a_n1186_n1046.n42 a_n1186_n1046.n41 2.7564
R501 a_n1186_n1046.n22 a_n1186_n1046.n10 2.64389
R502 a_n1186_n1046.n40 a_n1186_n1046.n34 2.13493
R503 a_n1186_n1046.n43 a_n1186_n1046.n40 1.60663
R504 a_n1186_n1046.n39 a_n1186_n1046.n38 1.04597
R505 a_n1186_n1046.n46 a_n1186_n1046.n45 0.802904
R506 a_n1186_n1046.n22 a_n1186_n1046.n21 0.768
R507 a_n1186_n1046.n33 a_n1186_n1046.n32 0.726409
R508 a_n1186_n1046.n38 a_n1186_n1046.n37 0.716442
R509 a_n1186_n1046.n36 a_n1186_n1046.n35 0.686026
R510 a_n1186_n1046.n49 a_n1186_n1046.n48 0.6155
R511 a_n1186_n1046.n29 a_n1186_n1046.n28 0.526182
R512 a_n1186_n1046.n30 a_n1186_n1046.n29 0.526182
R513 a_n1186_n1046.n31 a_n1186_n1046.n30 0.526182
R514 a_n1186_n1046.n32 a_n1186_n1046.n31 0.526182
R515 a_n1186_n1046.n24 a_n1186_n1046.n23 0.502015
R516 a_n1186_n1046.n25 a_n1186_n1046.n24 0.502015
R517 a_n1186_n1046.n26 a_n1186_n1046.n25 0.502015
R518 a_n1186_n1046.n27 a_n1186_n1046.n26 0.502015
R519 a_n1186_n1046.n21 a_n1186_n1046.n20 0.4805
R520 a_n1186_n1046.n20 a_n1186_n1046.n19 0.4805
R521 a_n1186_n1046.n19 a_n1186_n1046.n18 0.4805
R522 a_n1186_n1046.n18 a_n1186_n1046.n17 0.4805
R523 a_n1186_n1046.n17 a_n1186_n1046.n16 0.4805
R524 a_n1186_n1046.n16 a_n1186_n1046.n15 0.4805
R525 a_n1186_n1046.n15 a_n1186_n1046.n14 0.4805
R526 a_n1186_n1046.n14 a_n1186_n1046.n13 0.4805
R527 a_n1186_n1046.n13 a_n1186_n1046.n12 0.4805
R528 a_n1186_n1046.n12 a_n1186_n1046.n11 0.4805
R529 a_n1186_n1046.n1 a_n1186_n1046.n0 0.427272
R530 a_n1186_n1046.n2 a_n1186_n1046.n1 0.427272
R531 a_n1186_n1046.n3 a_n1186_n1046.n2 0.427272
R532 a_n1186_n1046.n4 a_n1186_n1046.n3 0.427272
R533 a_n1186_n1046.n5 a_n1186_n1046.n4 0.427272
R534 a_n1186_n1046.n6 a_n1186_n1046.n5 0.427272
R535 a_n1186_n1046.n7 a_n1186_n1046.n6 0.427272
R536 a_n1186_n1046.n8 a_n1186_n1046.n7 0.427272
R537 a_n1186_n1046.n9 a_n1186_n1046.n8 0.427272
R538 a_n1186_n1046.n10 a_n1186_n1046.n9 0.427272
R539 a_5585_876.n15 a_5585_876.t2 47.1257
R540 a_5585_876.n15 a_5585_876.n14 37.573
R541 a_5585_876.n1 a_5585_876.t7 36.1999
R542 a_5585_876.n16 a_5585_876.t11 31.1998
R543 a_5585_876.n18 a_5585_876.n17 29.4552
R544 a_5585_876.n24 a_5585_876.n23 29.4552
R545 a_5585_876.n22 a_5585_876.n21 29.4498
R546 a_5585_876.n20 a_5585_876.n19 29.4498
R547 a_5585_876.n13 a_5585_876.n12 29.4498
R548 a_5585_876.n11 a_5585_876.n10 29.4498
R549 a_5585_876.n9 a_5585_876.n8 29.4498
R550 a_5585_876.n7 a_5585_876.n6 29.4498
R551 a_5585_876.n5 a_5585_876.n4 29.4498
R552 a_5585_876.n3 a_5585_876.n2 29.4498
R553 a_5585_876.n1 a_5585_876.n0 29.4498
R554 a_5585_876.n16 a_5585_876.n15 11.4723
R555 a_5585_876.n14 a_5585_876.t0 9.0005
R556 a_5585_876.n14 a_5585_876.t1 9.0005
R557 a_5585_876.n21 a_5585_876.t9 6.2505
R558 a_5585_876.n21 a_5585_876.t12 6.2505
R559 a_5585_876.n19 a_5585_876.t13 6.2505
R560 a_5585_876.n19 a_5585_876.t23 6.2505
R561 a_5585_876.n17 a_5585_876.t26 6.2505
R562 a_5585_876.n17 a_5585_876.t4 6.2505
R563 a_5585_876.n12 a_5585_876.t17 6.2505
R564 a_5585_876.n12 a_5585_876.t20 6.2505
R565 a_5585_876.n10 a_5585_876.t6 6.2505
R566 a_5585_876.n10 a_5585_876.t14 6.2505
R567 a_5585_876.n8 a_5585_876.t24 6.2505
R568 a_5585_876.n8 a_5585_876.t5 6.2505
R569 a_5585_876.n6 a_5585_876.t16 6.2505
R570 a_5585_876.n6 a_5585_876.t19 6.2505
R571 a_5585_876.n4 a_5585_876.t3 6.2505
R572 a_5585_876.n4 a_5585_876.t10 6.2505
R573 a_5585_876.n2 a_5585_876.t18 6.2505
R574 a_5585_876.n2 a_5585_876.t22 6.2505
R575 a_5585_876.n0 a_5585_876.t8 6.2505
R576 a_5585_876.n0 a_5585_876.t15 6.2505
R577 a_5585_876.n24 a_5585_876.t21 6.2505
R578 a_5585_876.t25 a_5585_876.n24 6.2505
R579 a_5585_876.n18 a_5585_876.n16 4.99471
R580 a_5585_876.n20 a_5585_876.n18 0.506613
R581 a_5585_876.n23 a_5585_876.n22 0.494708
R582 a_5585_876.n3 a_5585_876.n1 0.494708
R583 a_5585_876.n5 a_5585_876.n3 0.494708
R584 a_5585_876.n9 a_5585_876.n7 0.494708
R585 a_5585_876.n11 a_5585_876.n9 0.494708
R586 a_5585_876.n13 a_5585_876.n11 0.494708
R587 a_5585_876.n23 a_5585_876.n13 0.494708
R588 a_5585_876.n22 a_5585_876.n20 0.488756
R589 a_5585_876.n7 a_5585_876.n5 0.488756
R590 D0.n1 D0.t2 483.342
R591 D0.n0 D0.t1 483.009
R592 D0.n0 D0.t0 482.634
R593 D0 D0.n1 2.38932
R594 D0.n1 D0.n0 1.43214
R595 D3.n1 D3.t2 483.75
R596 D3.n0 D3.t1 483.211
R597 D3.n0 D3.t0 482.634
R598 D3 D3.n1 5.76373
R599 D3.n1 D3.n0 2.28555
R600 Vref Vref.t0 43.0035
R601 VDD VDD.t0 22.553
R602 D1.n1 D1.t0 483.498
R603 D1.n0 D1.t2 483.034
R604 D1.n0 D1.t1 482.634
R605 D1 D1.n1 5.5923
R606 D1.n1 D1.n0 1.64842
C0 OUT VDD 0.024599f
C1 D2 a_3992_n1502# 0.311866f
C2 a_3992_n1502# a_2756_n1382# 0.033313f
C3 D1 a_3992_n1502# 0.020844f
C4 D2 OUT 0.561004f
C5 OUT a_2756_n1382# 1.07527f
C6 D1 OUT 0.54461f
C7 a_1632_n1418# OUT 1.08973f
C8 D3 a_3992_n1502# 1.76e-19
C9 D2 a_2756_n1382# 2.87e-20
C10 D2 D1 0.029366f
C11 D1 a_2756_n1382# 0.313829f
C12 D3 OUT 0.501139f
C13 a_1632_n1418# a_2756_n1382# 0.037834f
C14 D1 a_1632_n1418# 9.59e-20
C15 D2 D3 0.028012f
C16 D0 OUT 0.557993f
C17 D0 a_2756_n1382# 0.021996f
C18 D0 D1 0.033483f
C19 D0 a_1632_n1418# 0.342438f
C20 OUT a_3992_n1502# 1.08752f
C21 D3 VSS 1.53651f
C22 D2 VSS 1.49945f
C23 D1 VSS 1.58889f
C24 D0 VSS 1.71254f
C25 VDD VSS 1.29816f
C26 OUT VSS 4.78232f
C27 Vref VSS 0.98457f
C28 a_3992_n1502# VSS 7.53222f
C29 a_2756_n1382# VSS 4.48361f
C30 a_1632_n1418# VSS 2.99463f
C31 a_n1774_2554# VSS 1.49828f
C32 a_5585_876.t21 VSS 0.014204f
C33 a_5585_876.t7 VSS 0.061871f
C34 a_5585_876.t8 VSS 0.014204f
C35 a_5585_876.t15 VSS 0.014204f
C36 a_5585_876.n0 VSS 0.043095f
C37 a_5585_876.n1 VSS 0.164347f
C38 a_5585_876.t18 VSS 0.014204f
C39 a_5585_876.t22 VSS 0.014204f
C40 a_5585_876.n2 VSS 0.043095f
C41 a_5585_876.n3 VSS 0.08004f
C42 a_5585_876.t3 VSS 0.014204f
C43 a_5585_876.t10 VSS 0.014204f
C44 a_5585_876.n4 VSS 0.043095f
C45 a_5585_876.n5 VSS 0.079971f
C46 a_5585_876.t16 VSS 0.014204f
C47 a_5585_876.t19 VSS 0.014204f
C48 a_5585_876.n6 VSS 0.043095f
C49 a_5585_876.n7 VSS 0.079971f
C50 a_5585_876.t24 VSS 0.014204f
C51 a_5585_876.t5 VSS 0.014204f
C52 a_5585_876.n8 VSS 0.043095f
C53 a_5585_876.n9 VSS 0.08004f
C54 a_5585_876.t6 VSS 0.014204f
C55 a_5585_876.t14 VSS 0.014204f
C56 a_5585_876.n10 VSS 0.043095f
C57 a_5585_876.n11 VSS 0.08004f
C58 a_5585_876.t17 VSS 0.014204f
C59 a_5585_876.t20 VSS 0.014204f
C60 a_5585_876.n12 VSS 0.043095f
C61 a_5585_876.n13 VSS 0.08004f
C62 a_5585_876.t2 VSS 0.040307f
C63 a_5585_876.t0 VSS 0.009864f
C64 a_5585_876.t1 VSS 0.009864f
C65 a_5585_876.n14 VSS 0.027612f
C66 a_5585_876.n15 VSS 0.200666f
C67 a_5585_876.t11 VSS 0.050091f
C68 a_5585_876.n16 VSS 0.239262f
C69 a_5585_876.t26 VSS 0.014204f
C70 a_5585_876.t4 VSS 0.014204f
C71 a_5585_876.n17 VSS 0.043152f
C72 a_5585_876.n18 VSS 0.088992f
C73 a_5585_876.t13 VSS 0.014204f
C74 a_5585_876.t23 VSS 0.014204f
C75 a_5585_876.n19 VSS 0.043095f
C76 a_5585_876.n20 VSS 0.080109f
C77 a_5585_876.t9 VSS 0.014204f
C78 a_5585_876.t12 VSS 0.014204f
C79 a_5585_876.n21 VSS 0.043095f
C80 a_5585_876.n22 VSS 0.079971f
C81 a_5585_876.n23 VSS 0.080286f
C82 a_5585_876.n24 VSS 0.043152f
C83 a_5585_876.t25 VSS 0.014204f
C84 a_n1186_n1046.t37 VSS 0.01341f
C85 a_n1186_n1046.t9 VSS 0.013402f
C86 a_n1186_n1046.n0 VSS 0.026653f
C87 a_n1186_n1046.t34 VSS 0.013402f
C88 a_n1186_n1046.n1 VSS 0.015268f
C89 a_n1186_n1046.t39 VSS 0.013402f
C90 a_n1186_n1046.n2 VSS 0.015268f
C91 a_n1186_n1046.t16 VSS 0.013402f
C92 a_n1186_n1046.n3 VSS 0.015268f
C93 a_n1186_n1046.t23 VSS 0.013402f
C94 a_n1186_n1046.n4 VSS 0.015268f
C95 a_n1186_n1046.t43 VSS 0.013402f
C96 a_n1186_n1046.n5 VSS 0.015268f
C97 a_n1186_n1046.t11 VSS 0.013402f
C98 a_n1186_n1046.n6 VSS 0.015268f
C99 a_n1186_n1046.t24 VSS 0.013402f
C100 a_n1186_n1046.n7 VSS 0.015268f
C101 a_n1186_n1046.t48 VSS 0.013402f
C102 a_n1186_n1046.n8 VSS 0.015268f
C103 a_n1186_n1046.t20 VSS 0.013402f
C104 a_n1186_n1046.n9 VSS 0.015268f
C105 a_n1186_n1046.t40 VSS 0.013402f
C106 a_n1186_n1046.n10 VSS 0.032364f
C107 a_n1186_n1046.t47 VSS 0.013412f
C108 a_n1186_n1046.t14 VSS 0.013402f
C109 a_n1186_n1046.n11 VSS 0.027165f
C110 a_n1186_n1046.t35 VSS 0.013402f
C111 a_n1186_n1046.n12 VSS 0.014016f
C112 a_n1186_n1046.t10 VSS 0.013402f
C113 a_n1186_n1046.n13 VSS 0.014016f
C114 a_n1186_n1046.t17 VSS 0.013402f
C115 a_n1186_n1046.n14 VSS 0.014016f
C116 a_n1186_n1046.t30 VSS 0.013402f
C117 a_n1186_n1046.n15 VSS 0.014016f
C118 a_n1186_n1046.t44 VSS 0.013402f
C119 a_n1186_n1046.n16 VSS 0.014016f
C120 a_n1186_n1046.t18 VSS 0.013402f
C121 a_n1186_n1046.n17 VSS 0.014016f
C122 a_n1186_n1046.t38 VSS 0.013402f
C123 a_n1186_n1046.n18 VSS 0.014016f
C124 a_n1186_n1046.t15 VSS 0.013402f
C125 a_n1186_n1046.n19 VSS 0.014016f
C126 a_n1186_n1046.t26 VSS 0.013402f
C127 a_n1186_n1046.n20 VSS 0.014016f
C128 a_n1186_n1046.t41 VSS 0.013402f
C129 a_n1186_n1046.n21 VSS 0.016159f
C130 a_n1186_n1046.n22 VSS 0.093228f
C131 a_n1186_n1046.t31 VSS 0.012897f
C132 a_n1186_n1046.t50 VSS 0.012889f
C133 a_n1186_n1046.n23 VSS 0.023156f
C134 a_n1186_n1046.t25 VSS 0.012889f
C135 a_n1186_n1046.n24 VSS 0.013664f
C136 a_n1186_n1046.t49 VSS 0.012889f
C137 a_n1186_n1046.n25 VSS 0.013664f
C138 a_n1186_n1046.t22 VSS 0.012889f
C139 a_n1186_n1046.n26 VSS 0.013664f
C140 a_n1186_n1046.t29 VSS 0.012889f
C141 a_n1186_n1046.n27 VSS 0.027418f
C142 a_n1186_n1046.t46 VSS 0.012895f
C143 a_n1186_n1046.t19 VSS 0.012889f
C144 a_n1186_n1046.n28 VSS 0.019933f
C145 a_n1186_n1046.t32 VSS 0.012889f
C146 a_n1186_n1046.n29 VSS 0.013232f
C147 a_n1186_n1046.t51 VSS 0.012889f
C148 a_n1186_n1046.n30 VSS 0.013232f
C149 a_n1186_n1046.t28 VSS 0.012889f
C150 a_n1186_n1046.n31 VSS 0.013232f
C151 a_n1186_n1046.t42 VSS 0.012889f
C152 a_n1186_n1046.n32 VSS 0.014375f
C153 a_n1186_n1046.n33 VSS 0.038222f
C154 a_n1186_n1046.n34 VSS 0.268924f
C155 a_n1186_n1046.t36 VSS 0.012586f
C156 a_n1186_n1046.t8 VSS 0.012574f
C157 a_n1186_n1046.n35 VSS 0.022197f
C158 a_n1186_n1046.t13 VSS 0.012574f
C159 a_n1186_n1046.n36 VSS 0.021373f
C160 a_n1186_n1046.t45 VSS 0.012583f
C161 a_n1186_n1046.t12 VSS 0.012574f
C162 a_n1186_n1046.n37 VSS 0.018368f
C163 a_n1186_n1046.t21 VSS 0.012574f
C164 a_n1186_n1046.n38 VSS 0.01241f
C165 a_n1186_n1046.n39 VSS 0.024502f
C166 a_n1186_n1046.n40 VSS 0.127329f
C167 a_n1186_n1046.t7 VSS 0.012582f
C168 a_n1186_n1046.t33 VSS 0.012574f
C169 a_n1186_n1046.n41 VSS 0.033248f
C170 a_n1186_n1046.t27 VSS 0.012594f
C171 a_n1186_n1046.n42 VSS 0.04594f
C172 a_n1186_n1046.n43 VSS 0.145194f
C173 a_n1186_n1046.t4 VSS 0.012586f
C174 a_n1186_n1046.t0 VSS 0.012574f
C175 a_n1186_n1046.n44 VSS 0.02823f
C176 a_n1186_n1046.t2 VSS 0.012597f
C177 a_n1186_n1046.n45 VSS 0.027952f
C178 a_n1186_n1046.n46 VSS 0.085967f
C179 a_n1186_n1046.t1 VSS 0.005969f
C180 a_n1186_n1046.t3 VSS 0.005969f
C181 a_n1186_n1046.n47 VSS 0.023491f
C182 a_n1186_n1046.t5 VSS 0.020832f
C183 a_n1186_n1046.n48 VSS 0.072068f
C184 a_n1186_n1046.n49 VSS 0.064608f
C185 a_n1186_n1046.t6 VSS 0.055192f
.ends
.end
