magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -631 -560 631 560
<< nmos >>
rect -445 -422 -345 360
rect -287 -422 -187 360
rect -129 -422 -29 360
rect 29 -422 129 360
rect 187 -422 287 360
rect 345 -422 445 360
<< ndiff >>
rect -503 326 -445 360
rect -503 292 -491 326
rect -457 292 -445 326
rect -503 258 -445 292
rect -503 224 -491 258
rect -457 224 -445 258
rect -503 190 -445 224
rect -503 156 -491 190
rect -457 156 -445 190
rect -503 122 -445 156
rect -503 88 -491 122
rect -457 88 -445 122
rect -503 54 -445 88
rect -503 20 -491 54
rect -457 20 -445 54
rect -503 -14 -445 20
rect -503 -48 -491 -14
rect -457 -48 -445 -14
rect -503 -82 -445 -48
rect -503 -116 -491 -82
rect -457 -116 -445 -82
rect -503 -150 -445 -116
rect -503 -184 -491 -150
rect -457 -184 -445 -150
rect -503 -218 -445 -184
rect -503 -252 -491 -218
rect -457 -252 -445 -218
rect -503 -286 -445 -252
rect -503 -320 -491 -286
rect -457 -320 -445 -286
rect -503 -354 -445 -320
rect -503 -388 -491 -354
rect -457 -388 -445 -354
rect -503 -422 -445 -388
rect -345 326 -287 360
rect -345 292 -333 326
rect -299 292 -287 326
rect -345 258 -287 292
rect -345 224 -333 258
rect -299 224 -287 258
rect -345 190 -287 224
rect -345 156 -333 190
rect -299 156 -287 190
rect -345 122 -287 156
rect -345 88 -333 122
rect -299 88 -287 122
rect -345 54 -287 88
rect -345 20 -333 54
rect -299 20 -287 54
rect -345 -14 -287 20
rect -345 -48 -333 -14
rect -299 -48 -287 -14
rect -345 -82 -287 -48
rect -345 -116 -333 -82
rect -299 -116 -287 -82
rect -345 -150 -287 -116
rect -345 -184 -333 -150
rect -299 -184 -287 -150
rect -345 -218 -287 -184
rect -345 -252 -333 -218
rect -299 -252 -287 -218
rect -345 -286 -287 -252
rect -345 -320 -333 -286
rect -299 -320 -287 -286
rect -345 -354 -287 -320
rect -345 -388 -333 -354
rect -299 -388 -287 -354
rect -345 -422 -287 -388
rect -187 326 -129 360
rect -187 292 -175 326
rect -141 292 -129 326
rect -187 258 -129 292
rect -187 224 -175 258
rect -141 224 -129 258
rect -187 190 -129 224
rect -187 156 -175 190
rect -141 156 -129 190
rect -187 122 -129 156
rect -187 88 -175 122
rect -141 88 -129 122
rect -187 54 -129 88
rect -187 20 -175 54
rect -141 20 -129 54
rect -187 -14 -129 20
rect -187 -48 -175 -14
rect -141 -48 -129 -14
rect -187 -82 -129 -48
rect -187 -116 -175 -82
rect -141 -116 -129 -82
rect -187 -150 -129 -116
rect -187 -184 -175 -150
rect -141 -184 -129 -150
rect -187 -218 -129 -184
rect -187 -252 -175 -218
rect -141 -252 -129 -218
rect -187 -286 -129 -252
rect -187 -320 -175 -286
rect -141 -320 -129 -286
rect -187 -354 -129 -320
rect -187 -388 -175 -354
rect -141 -388 -129 -354
rect -187 -422 -129 -388
rect -29 326 29 360
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -422 29 -388
rect 129 326 187 360
rect 129 292 141 326
rect 175 292 187 326
rect 129 258 187 292
rect 129 224 141 258
rect 175 224 187 258
rect 129 190 187 224
rect 129 156 141 190
rect 175 156 187 190
rect 129 122 187 156
rect 129 88 141 122
rect 175 88 187 122
rect 129 54 187 88
rect 129 20 141 54
rect 175 20 187 54
rect 129 -14 187 20
rect 129 -48 141 -14
rect 175 -48 187 -14
rect 129 -82 187 -48
rect 129 -116 141 -82
rect 175 -116 187 -82
rect 129 -150 187 -116
rect 129 -184 141 -150
rect 175 -184 187 -150
rect 129 -218 187 -184
rect 129 -252 141 -218
rect 175 -252 187 -218
rect 129 -286 187 -252
rect 129 -320 141 -286
rect 175 -320 187 -286
rect 129 -354 187 -320
rect 129 -388 141 -354
rect 175 -388 187 -354
rect 129 -422 187 -388
rect 287 326 345 360
rect 287 292 299 326
rect 333 292 345 326
rect 287 258 345 292
rect 287 224 299 258
rect 333 224 345 258
rect 287 190 345 224
rect 287 156 299 190
rect 333 156 345 190
rect 287 122 345 156
rect 287 88 299 122
rect 333 88 345 122
rect 287 54 345 88
rect 287 20 299 54
rect 333 20 345 54
rect 287 -14 345 20
rect 287 -48 299 -14
rect 333 -48 345 -14
rect 287 -82 345 -48
rect 287 -116 299 -82
rect 333 -116 345 -82
rect 287 -150 345 -116
rect 287 -184 299 -150
rect 333 -184 345 -150
rect 287 -218 345 -184
rect 287 -252 299 -218
rect 333 -252 345 -218
rect 287 -286 345 -252
rect 287 -320 299 -286
rect 333 -320 345 -286
rect 287 -354 345 -320
rect 287 -388 299 -354
rect 333 -388 345 -354
rect 287 -422 345 -388
rect 445 326 503 360
rect 445 292 457 326
rect 491 292 503 326
rect 445 258 503 292
rect 445 224 457 258
rect 491 224 503 258
rect 445 190 503 224
rect 445 156 457 190
rect 491 156 503 190
rect 445 122 503 156
rect 445 88 457 122
rect 491 88 503 122
rect 445 54 503 88
rect 445 20 457 54
rect 491 20 503 54
rect 445 -14 503 20
rect 445 -48 457 -14
rect 491 -48 503 -14
rect 445 -82 503 -48
rect 445 -116 457 -82
rect 491 -116 503 -82
rect 445 -150 503 -116
rect 445 -184 457 -150
rect 491 -184 503 -150
rect 445 -218 503 -184
rect 445 -252 457 -218
rect 491 -252 503 -218
rect 445 -286 503 -252
rect 445 -320 457 -286
rect 491 -320 503 -286
rect 445 -354 503 -320
rect 445 -388 457 -354
rect 491 -388 503 -354
rect 445 -422 503 -388
<< ndiffc >>
rect -491 292 -457 326
rect -491 224 -457 258
rect -491 156 -457 190
rect -491 88 -457 122
rect -491 20 -457 54
rect -491 -48 -457 -14
rect -491 -116 -457 -82
rect -491 -184 -457 -150
rect -491 -252 -457 -218
rect -491 -320 -457 -286
rect -491 -388 -457 -354
rect -333 292 -299 326
rect -333 224 -299 258
rect -333 156 -299 190
rect -333 88 -299 122
rect -333 20 -299 54
rect -333 -48 -299 -14
rect -333 -116 -299 -82
rect -333 -184 -299 -150
rect -333 -252 -299 -218
rect -333 -320 -299 -286
rect -333 -388 -299 -354
rect -175 292 -141 326
rect -175 224 -141 258
rect -175 156 -141 190
rect -175 88 -141 122
rect -175 20 -141 54
rect -175 -48 -141 -14
rect -175 -116 -141 -82
rect -175 -184 -141 -150
rect -175 -252 -141 -218
rect -175 -320 -141 -286
rect -175 -388 -141 -354
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect 141 292 175 326
rect 141 224 175 258
rect 141 156 175 190
rect 141 88 175 122
rect 141 20 175 54
rect 141 -48 175 -14
rect 141 -116 175 -82
rect 141 -184 175 -150
rect 141 -252 175 -218
rect 141 -320 175 -286
rect 141 -388 175 -354
rect 299 292 333 326
rect 299 224 333 258
rect 299 156 333 190
rect 299 88 333 122
rect 299 20 333 54
rect 299 -48 333 -14
rect 299 -116 333 -82
rect 299 -184 333 -150
rect 299 -252 333 -218
rect 299 -320 333 -286
rect 299 -388 333 -354
rect 457 292 491 326
rect 457 224 491 258
rect 457 156 491 190
rect 457 88 491 122
rect 457 20 491 54
rect 457 -48 491 -14
rect 457 -116 491 -82
rect 457 -184 491 -150
rect 457 -252 491 -218
rect 457 -320 491 -286
rect 457 -388 491 -354
<< psubdiff >>
rect -605 500 -493 534
rect -459 500 -425 534
rect -391 500 -357 534
rect -323 500 -289 534
rect -255 500 -221 534
rect -187 500 -153 534
rect -119 500 -85 534
rect -51 500 -17 534
rect 17 500 51 534
rect 85 500 119 534
rect 153 500 187 534
rect 221 500 255 534
rect 289 500 323 534
rect 357 500 391 534
rect 425 500 459 534
rect 493 500 605 534
rect -605 425 -571 500
rect -605 357 -571 391
rect 571 425 605 500
rect -605 289 -571 323
rect -605 221 -571 255
rect -605 153 -571 187
rect -605 85 -571 119
rect -605 17 -571 51
rect -605 -51 -571 -17
rect -605 -119 -571 -85
rect -605 -187 -571 -153
rect -605 -255 -571 -221
rect -605 -323 -571 -289
rect -605 -391 -571 -357
rect 571 357 605 391
rect 571 289 605 323
rect 571 221 605 255
rect 571 153 605 187
rect 571 85 605 119
rect 571 17 605 51
rect 571 -51 605 -17
rect 571 -119 605 -85
rect 571 -187 605 -153
rect 571 -255 605 -221
rect 571 -323 605 -289
rect 571 -391 605 -357
rect -605 -500 -571 -425
rect 571 -500 605 -425
rect -605 -534 -493 -500
rect -459 -534 -425 -500
rect -391 -534 -357 -500
rect -323 -534 -289 -500
rect -255 -534 -221 -500
rect -187 -534 -153 -500
rect -119 -534 -85 -500
rect -51 -534 -17 -500
rect 17 -534 51 -500
rect 85 -534 119 -500
rect 153 -534 187 -500
rect 221 -534 255 -500
rect 289 -534 323 -500
rect 357 -534 391 -500
rect 425 -534 459 -500
rect 493 -534 605 -500
<< psubdiffcont >>
rect -493 500 -459 534
rect -425 500 -391 534
rect -357 500 -323 534
rect -289 500 -255 534
rect -221 500 -187 534
rect -153 500 -119 534
rect -85 500 -51 534
rect -17 500 17 534
rect 51 500 85 534
rect 119 500 153 534
rect 187 500 221 534
rect 255 500 289 534
rect 323 500 357 534
rect 391 500 425 534
rect 459 500 493 534
rect -605 391 -571 425
rect 571 391 605 425
rect -605 323 -571 357
rect -605 255 -571 289
rect -605 187 -571 221
rect -605 119 -571 153
rect -605 51 -571 85
rect -605 -17 -571 17
rect -605 -85 -571 -51
rect -605 -153 -571 -119
rect -605 -221 -571 -187
rect -605 -289 -571 -255
rect -605 -357 -571 -323
rect -605 -425 -571 -391
rect 571 323 605 357
rect 571 255 605 289
rect 571 187 605 221
rect 571 119 605 153
rect 571 51 605 85
rect 571 -17 605 17
rect 571 -85 605 -51
rect 571 -153 605 -119
rect 571 -221 605 -187
rect 571 -289 605 -255
rect 571 -357 605 -323
rect 571 -425 605 -391
rect -493 -534 -459 -500
rect -425 -534 -391 -500
rect -357 -534 -323 -500
rect -289 -534 -255 -500
rect -221 -534 -187 -500
rect -153 -534 -119 -500
rect -85 -534 -51 -500
rect -17 -534 17 -500
rect 51 -534 85 -500
rect 119 -534 153 -500
rect 187 -534 221 -500
rect 255 -534 289 -500
rect 323 -534 357 -500
rect 391 -534 425 -500
rect 459 -534 493 -500
<< poly >>
rect -445 432 -345 448
rect -445 398 -412 432
rect -378 398 -345 432
rect -445 360 -345 398
rect -287 432 -187 448
rect -287 398 -254 432
rect -220 398 -187 432
rect -287 360 -187 398
rect -129 432 -29 448
rect -129 398 -96 432
rect -62 398 -29 432
rect -129 360 -29 398
rect 29 432 129 448
rect 29 398 62 432
rect 96 398 129 432
rect 29 360 129 398
rect 187 432 287 448
rect 187 398 220 432
rect 254 398 287 432
rect 187 360 287 398
rect 345 432 445 448
rect 345 398 378 432
rect 412 398 445 432
rect 345 360 445 398
rect -445 -448 -345 -422
rect -287 -448 -187 -422
rect -129 -448 -29 -422
rect 29 -448 129 -422
rect 187 -448 287 -422
rect 345 -448 445 -422
<< polycont >>
rect -412 398 -378 432
rect -254 398 -220 432
rect -96 398 -62 432
rect 62 398 96 432
rect 220 398 254 432
rect 378 398 412 432
<< locali >>
rect -605 500 -493 534
rect -459 500 -425 534
rect -391 500 -357 534
rect -323 500 -289 534
rect -255 500 -221 534
rect -187 500 -153 534
rect -119 500 -85 534
rect -51 500 -17 534
rect 17 500 51 534
rect 85 500 119 534
rect 153 500 187 534
rect 221 500 255 534
rect 289 500 323 534
rect 357 500 391 534
rect 425 500 459 534
rect 493 500 605 534
rect -605 425 -571 500
rect -445 398 -412 432
rect -378 398 -345 432
rect -287 398 -254 432
rect -220 398 -187 432
rect -129 398 -96 432
rect -62 398 -29 432
rect 29 398 62 432
rect 96 398 129 432
rect 187 398 220 432
rect 254 398 287 432
rect 345 398 378 432
rect 412 398 445 432
rect 571 425 605 500
rect -605 357 -571 391
rect -605 289 -571 323
rect -605 221 -571 255
rect -605 153 -571 187
rect -605 85 -571 119
rect -605 17 -571 51
rect -605 -51 -571 -17
rect -605 -119 -571 -85
rect -605 -187 -571 -153
rect -605 -255 -571 -221
rect -605 -323 -571 -289
rect -605 -391 -571 -357
rect -605 -500 -571 -425
rect -491 346 -457 364
rect -491 274 -457 292
rect -491 202 -457 224
rect -491 130 -457 156
rect -491 58 -457 88
rect -491 -14 -457 20
rect -491 -82 -457 -48
rect -491 -150 -457 -120
rect -491 -218 -457 -192
rect -491 -286 -457 -264
rect -491 -354 -457 -336
rect -491 -426 -457 -408
rect -333 346 -299 364
rect -333 274 -299 292
rect -333 202 -299 224
rect -333 130 -299 156
rect -333 58 -299 88
rect -333 -14 -299 20
rect -333 -82 -299 -48
rect -333 -150 -299 -120
rect -333 -218 -299 -192
rect -333 -286 -299 -264
rect -333 -354 -299 -336
rect -333 -426 -299 -408
rect -175 346 -141 364
rect -175 274 -141 292
rect -175 202 -141 224
rect -175 130 -141 156
rect -175 58 -141 88
rect -175 -14 -141 20
rect -175 -82 -141 -48
rect -175 -150 -141 -120
rect -175 -218 -141 -192
rect -175 -286 -141 -264
rect -175 -354 -141 -336
rect -175 -426 -141 -408
rect -17 346 17 364
rect -17 274 17 292
rect -17 202 17 224
rect -17 130 17 156
rect -17 58 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -120
rect -17 -218 17 -192
rect -17 -286 17 -264
rect -17 -354 17 -336
rect -17 -426 17 -408
rect 141 346 175 364
rect 141 274 175 292
rect 141 202 175 224
rect 141 130 175 156
rect 141 58 175 88
rect 141 -14 175 20
rect 141 -82 175 -48
rect 141 -150 175 -120
rect 141 -218 175 -192
rect 141 -286 175 -264
rect 141 -354 175 -336
rect 141 -426 175 -408
rect 299 346 333 364
rect 299 274 333 292
rect 299 202 333 224
rect 299 130 333 156
rect 299 58 333 88
rect 299 -14 333 20
rect 299 -82 333 -48
rect 299 -150 333 -120
rect 299 -218 333 -192
rect 299 -286 333 -264
rect 299 -354 333 -336
rect 299 -426 333 -408
rect 457 346 491 364
rect 457 274 491 292
rect 457 202 491 224
rect 457 130 491 156
rect 457 58 491 88
rect 457 -14 491 20
rect 457 -82 491 -48
rect 457 -150 491 -120
rect 457 -218 491 -192
rect 457 -286 491 -264
rect 457 -354 491 -336
rect 457 -426 491 -408
rect 571 357 605 391
rect 571 289 605 323
rect 571 221 605 255
rect 571 153 605 187
rect 571 85 605 119
rect 571 17 605 51
rect 571 -51 605 -17
rect 571 -119 605 -85
rect 571 -187 605 -153
rect 571 -255 605 -221
rect 571 -323 605 -289
rect 571 -391 605 -357
rect 571 -500 605 -425
rect -605 -534 -493 -500
rect -459 -534 -425 -500
rect -391 -534 -357 -500
rect -323 -534 -289 -500
rect -255 -534 -221 -500
rect -187 -534 -153 -500
rect -119 -534 -85 -500
rect -51 -534 -17 -500
rect 17 -534 51 -500
rect 85 -534 119 -500
rect 153 -534 187 -500
rect 221 -534 255 -500
rect 289 -534 323 -500
rect 357 -534 391 -500
rect 425 -534 459 -500
rect 493 -534 605 -500
<< viali >>
rect -412 398 -378 432
rect -254 398 -220 432
rect -96 398 -62 432
rect 62 398 96 432
rect 220 398 254 432
rect 378 398 412 432
rect -491 326 -457 346
rect -491 312 -457 326
rect -491 258 -457 274
rect -491 240 -457 258
rect -491 190 -457 202
rect -491 168 -457 190
rect -491 122 -457 130
rect -491 96 -457 122
rect -491 54 -457 58
rect -491 24 -457 54
rect -491 -48 -457 -14
rect -491 -116 -457 -86
rect -491 -120 -457 -116
rect -491 -184 -457 -158
rect -491 -192 -457 -184
rect -491 -252 -457 -230
rect -491 -264 -457 -252
rect -491 -320 -457 -302
rect -491 -336 -457 -320
rect -491 -388 -457 -374
rect -491 -408 -457 -388
rect -333 326 -299 346
rect -333 312 -299 326
rect -333 258 -299 274
rect -333 240 -299 258
rect -333 190 -299 202
rect -333 168 -299 190
rect -333 122 -299 130
rect -333 96 -299 122
rect -333 54 -299 58
rect -333 24 -299 54
rect -333 -48 -299 -14
rect -333 -116 -299 -86
rect -333 -120 -299 -116
rect -333 -184 -299 -158
rect -333 -192 -299 -184
rect -333 -252 -299 -230
rect -333 -264 -299 -252
rect -333 -320 -299 -302
rect -333 -336 -299 -320
rect -333 -388 -299 -374
rect -333 -408 -299 -388
rect -175 326 -141 346
rect -175 312 -141 326
rect -175 258 -141 274
rect -175 240 -141 258
rect -175 190 -141 202
rect -175 168 -141 190
rect -175 122 -141 130
rect -175 96 -141 122
rect -175 54 -141 58
rect -175 24 -141 54
rect -175 -48 -141 -14
rect -175 -116 -141 -86
rect -175 -120 -141 -116
rect -175 -184 -141 -158
rect -175 -192 -141 -184
rect -175 -252 -141 -230
rect -175 -264 -141 -252
rect -175 -320 -141 -302
rect -175 -336 -141 -320
rect -175 -388 -141 -374
rect -175 -408 -141 -388
rect -17 326 17 346
rect -17 312 17 326
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect -17 -388 17 -374
rect -17 -408 17 -388
rect 141 326 175 346
rect 141 312 175 326
rect 141 258 175 274
rect 141 240 175 258
rect 141 190 175 202
rect 141 168 175 190
rect 141 122 175 130
rect 141 96 175 122
rect 141 54 175 58
rect 141 24 175 54
rect 141 -48 175 -14
rect 141 -116 175 -86
rect 141 -120 175 -116
rect 141 -184 175 -158
rect 141 -192 175 -184
rect 141 -252 175 -230
rect 141 -264 175 -252
rect 141 -320 175 -302
rect 141 -336 175 -320
rect 141 -388 175 -374
rect 141 -408 175 -388
rect 299 326 333 346
rect 299 312 333 326
rect 299 258 333 274
rect 299 240 333 258
rect 299 190 333 202
rect 299 168 333 190
rect 299 122 333 130
rect 299 96 333 122
rect 299 54 333 58
rect 299 24 333 54
rect 299 -48 333 -14
rect 299 -116 333 -86
rect 299 -120 333 -116
rect 299 -184 333 -158
rect 299 -192 333 -184
rect 299 -252 333 -230
rect 299 -264 333 -252
rect 299 -320 333 -302
rect 299 -336 333 -320
rect 299 -388 333 -374
rect 299 -408 333 -388
rect 457 326 491 346
rect 457 312 491 326
rect 457 258 491 274
rect 457 240 491 258
rect 457 190 491 202
rect 457 168 491 190
rect 457 122 491 130
rect 457 96 491 122
rect 457 54 491 58
rect 457 24 491 54
rect 457 -48 491 -14
rect 457 -116 491 -86
rect 457 -120 491 -116
rect 457 -184 491 -158
rect 457 -192 491 -184
rect 457 -252 491 -230
rect 457 -264 491 -252
rect 457 -320 491 -302
rect 457 -336 491 -320
rect 457 -388 491 -374
rect 457 -408 491 -388
<< metal1 >>
rect -441 432 -349 438
rect -441 398 -412 432
rect -378 398 -349 432
rect -441 392 -349 398
rect -283 432 -191 438
rect -283 398 -254 432
rect -220 398 -191 432
rect -283 392 -191 398
rect -125 432 -33 438
rect -125 398 -96 432
rect -62 398 -33 432
rect -125 392 -33 398
rect 33 432 125 438
rect 33 398 62 432
rect 96 398 125 432
rect 33 392 125 398
rect 191 432 283 438
rect 191 398 220 432
rect 254 398 283 432
rect 191 392 283 398
rect 349 432 441 438
rect 349 398 378 432
rect 412 398 441 432
rect 349 392 441 398
rect -497 346 -451 360
rect -497 312 -491 346
rect -457 312 -451 346
rect -497 274 -451 312
rect -497 240 -491 274
rect -457 240 -451 274
rect -497 202 -451 240
rect -497 168 -491 202
rect -457 168 -451 202
rect -497 130 -451 168
rect -497 96 -491 130
rect -457 96 -451 130
rect -497 58 -451 96
rect -497 24 -491 58
rect -457 24 -451 58
rect -497 -14 -451 24
rect -497 -48 -491 -14
rect -457 -48 -451 -14
rect -497 -86 -451 -48
rect -497 -120 -491 -86
rect -457 -120 -451 -86
rect -497 -158 -451 -120
rect -497 -192 -491 -158
rect -457 -192 -451 -158
rect -497 -230 -451 -192
rect -497 -264 -491 -230
rect -457 -264 -451 -230
rect -497 -302 -451 -264
rect -497 -336 -491 -302
rect -457 -336 -451 -302
rect -497 -374 -451 -336
rect -497 -408 -491 -374
rect -457 -408 -451 -374
rect -497 -422 -451 -408
rect -339 346 -293 360
rect -339 312 -333 346
rect -299 312 -293 346
rect -339 274 -293 312
rect -339 240 -333 274
rect -299 240 -293 274
rect -339 202 -293 240
rect -339 168 -333 202
rect -299 168 -293 202
rect -339 130 -293 168
rect -339 96 -333 130
rect -299 96 -293 130
rect -339 58 -293 96
rect -339 24 -333 58
rect -299 24 -293 58
rect -339 -14 -293 24
rect -339 -48 -333 -14
rect -299 -48 -293 -14
rect -339 -86 -293 -48
rect -339 -120 -333 -86
rect -299 -120 -293 -86
rect -339 -158 -293 -120
rect -339 -192 -333 -158
rect -299 -192 -293 -158
rect -339 -230 -293 -192
rect -339 -264 -333 -230
rect -299 -264 -293 -230
rect -339 -302 -293 -264
rect -339 -336 -333 -302
rect -299 -336 -293 -302
rect -339 -374 -293 -336
rect -339 -408 -333 -374
rect -299 -408 -293 -374
rect -339 -422 -293 -408
rect -181 346 -135 360
rect -181 312 -175 346
rect -141 312 -135 346
rect -181 274 -135 312
rect -181 240 -175 274
rect -141 240 -135 274
rect -181 202 -135 240
rect -181 168 -175 202
rect -141 168 -135 202
rect -181 130 -135 168
rect -181 96 -175 130
rect -141 96 -135 130
rect -181 58 -135 96
rect -181 24 -175 58
rect -141 24 -135 58
rect -181 -14 -135 24
rect -181 -48 -175 -14
rect -141 -48 -135 -14
rect -181 -86 -135 -48
rect -181 -120 -175 -86
rect -141 -120 -135 -86
rect -181 -158 -135 -120
rect -181 -192 -175 -158
rect -141 -192 -135 -158
rect -181 -230 -135 -192
rect -181 -264 -175 -230
rect -141 -264 -135 -230
rect -181 -302 -135 -264
rect -181 -336 -175 -302
rect -141 -336 -135 -302
rect -181 -374 -135 -336
rect -181 -408 -175 -374
rect -141 -408 -135 -374
rect -181 -422 -135 -408
rect -23 346 23 360
rect -23 312 -17 346
rect 17 312 23 346
rect -23 274 23 312
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -374 23 -336
rect -23 -408 -17 -374
rect 17 -408 23 -374
rect -23 -422 23 -408
rect 135 346 181 360
rect 135 312 141 346
rect 175 312 181 346
rect 135 274 181 312
rect 135 240 141 274
rect 175 240 181 274
rect 135 202 181 240
rect 135 168 141 202
rect 175 168 181 202
rect 135 130 181 168
rect 135 96 141 130
rect 175 96 181 130
rect 135 58 181 96
rect 135 24 141 58
rect 175 24 181 58
rect 135 -14 181 24
rect 135 -48 141 -14
rect 175 -48 181 -14
rect 135 -86 181 -48
rect 135 -120 141 -86
rect 175 -120 181 -86
rect 135 -158 181 -120
rect 135 -192 141 -158
rect 175 -192 181 -158
rect 135 -230 181 -192
rect 135 -264 141 -230
rect 175 -264 181 -230
rect 135 -302 181 -264
rect 135 -336 141 -302
rect 175 -336 181 -302
rect 135 -374 181 -336
rect 135 -408 141 -374
rect 175 -408 181 -374
rect 135 -422 181 -408
rect 293 346 339 360
rect 293 312 299 346
rect 333 312 339 346
rect 293 274 339 312
rect 293 240 299 274
rect 333 240 339 274
rect 293 202 339 240
rect 293 168 299 202
rect 333 168 339 202
rect 293 130 339 168
rect 293 96 299 130
rect 333 96 339 130
rect 293 58 339 96
rect 293 24 299 58
rect 333 24 339 58
rect 293 -14 339 24
rect 293 -48 299 -14
rect 333 -48 339 -14
rect 293 -86 339 -48
rect 293 -120 299 -86
rect 333 -120 339 -86
rect 293 -158 339 -120
rect 293 -192 299 -158
rect 333 -192 339 -158
rect 293 -230 339 -192
rect 293 -264 299 -230
rect 333 -264 339 -230
rect 293 -302 339 -264
rect 293 -336 299 -302
rect 333 -336 339 -302
rect 293 -374 339 -336
rect 293 -408 299 -374
rect 333 -408 339 -374
rect 293 -422 339 -408
rect 451 346 497 360
rect 451 312 457 346
rect 491 312 497 346
rect 451 274 497 312
rect 451 240 457 274
rect 491 240 497 274
rect 451 202 497 240
rect 451 168 457 202
rect 491 168 497 202
rect 451 130 497 168
rect 451 96 457 130
rect 491 96 497 130
rect 451 58 497 96
rect 451 24 457 58
rect 491 24 497 58
rect 451 -14 497 24
rect 451 -48 457 -14
rect 491 -48 497 -14
rect 451 -86 497 -48
rect 451 -120 457 -86
rect 491 -120 497 -86
rect 451 -158 497 -120
rect 451 -192 457 -158
rect 491 -192 497 -158
rect 451 -230 497 -192
rect 451 -264 457 -230
rect 491 -264 497 -230
rect 451 -302 497 -264
rect 451 -336 457 -302
rect 491 -336 497 -302
rect 451 -374 497 -336
rect 451 -408 457 -374
rect 491 -408 497 -374
rect 451 -422 497 -408
<< properties >>
string FIXED_BBOX -588 -517 588 517
<< end >>
