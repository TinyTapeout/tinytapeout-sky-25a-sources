magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -297 608 297 694
rect -297 -608 -211 608
rect 211 -608 297 608
rect -297 -694 297 -608
<< psubdiff >>
rect -271 634 -153 668
rect -119 634 -85 668
rect -51 634 -17 668
rect 17 634 51 668
rect 85 634 119 668
rect 153 634 271 668
rect -271 561 -237 634
rect 237 561 271 634
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect -271 -634 -237 -561
rect 237 -634 271 -561
rect -271 -668 -153 -634
rect -119 -668 -85 -634
rect -51 -668 -17 -634
rect 17 -668 51 -634
rect 85 -668 119 -634
rect 153 -668 271 -634
<< psubdiffcont >>
rect -153 634 -119 668
rect -85 634 -51 668
rect -17 634 17 668
rect 51 634 85 668
rect 119 634 153 668
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect -153 -668 -119 -634
rect -85 -668 -51 -634
rect -17 -668 17 -634
rect 51 -668 85 -634
rect 119 -668 153 -634
<< xpolycontact >>
rect -141 106 141 538
rect -141 -538 141 -106
<< xpolyres >>
rect -141 -106 141 106
<< locali >>
rect -271 634 -153 668
rect -119 634 -85 668
rect -51 634 -17 668
rect 17 634 51 668
rect 85 634 119 668
rect 153 634 271 668
rect -271 561 -237 634
rect 237 561 271 634
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect -271 -634 -237 -561
rect 237 -634 271 -561
rect -271 -668 -153 -634
rect -119 -668 -85 -634
rect -51 -668 -17 -634
rect 17 -668 51 -634
rect 85 -668 119 -634
rect 153 -668 271 -634
<< viali >>
rect -125 124 125 518
rect -125 -519 125 -125
<< metal1 >>
rect -131 518 131 532
rect -131 124 -125 518
rect 125 124 131 518
rect -131 111 131 124
rect -131 -125 131 -111
rect -131 -519 -125 -125
rect 125 -519 131 -125
rect -131 -532 131 -519
<< properties >>
string FIXED_BBOX -254 -651 254 651
<< end >>
