Incrementer Simulation
.include "pdk_lib.spice"

* instantiate the incrementer
*  
Xinc CLK VPWR RSTN INC VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND VGND OE0 OE1 OE2 OE3 OE4 OE5 OE6 OE7 S8 S9 S10 S11 S12 S13 S14 S15 S0 S1 S2 S3 S4 S5 S6 S7 VPWR VGND  tt_um_flat
