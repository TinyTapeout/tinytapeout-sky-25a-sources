magic
tech sky130A
timestamp 1757259598
<< metal4 >>
rect 6120 11160 6280 11320
rect 7160 11200 7280 11240
rect 7160 11160 7320 11200
rect 6120 11000 6320 11160
rect 7120 11120 7320 11160
rect 7120 11040 7360 11120
rect 6120 10880 6360 11000
rect 7080 10920 7400 11040
rect 6120 10760 6400 10880
rect 7080 10840 7440 10920
rect 6120 10720 6440 10760
rect 6160 10680 6440 10720
rect 7080 10680 7240 10840
rect 7280 10800 7480 10840
rect 7320 10760 7480 10800
rect 7320 10720 7520 10760
rect 7360 10680 7520 10720
rect 6160 10600 6480 10680
rect 6160 10520 6520 10600
rect 6200 10480 6560 10520
rect 6200 10360 6360 10480
rect 6400 10440 6600 10480
rect 7040 10440 7200 10680
rect 7360 10640 7560 10680
rect 7400 10600 7600 10640
rect 7440 10560 7600 10600
rect 7440 10520 7640 10560
rect 7480 10480 7680 10520
rect 7520 10440 7720 10480
rect 6440 10360 6640 10440
rect 6240 9600 6400 10360
rect 6480 10320 6680 10360
rect 6520 10240 6720 10320
rect 7000 10280 7160 10440
rect 7560 10400 7720 10440
rect 7560 10360 7760 10400
rect 7520 10320 7800 10360
rect 7440 10280 7840 10320
rect 6560 10200 6760 10240
rect 6600 10160 6800 10200
rect 6960 10160 7120 10280
rect 7360 10240 7880 10280
rect 7280 10200 7600 10240
rect 7680 10200 7920 10240
rect 7200 10160 7560 10200
rect 7720 10160 7960 10200
rect 6640 10120 6840 10160
rect 6920 10120 7120 10160
rect 7160 10120 7480 10160
rect 7760 10120 8000 10160
rect 6640 10080 6880 10120
rect 6920 10080 7080 10120
rect 6680 10040 7080 10080
rect 7160 10080 7400 10120
rect 7800 10080 8040 10120
rect 7160 10040 7320 10080
rect 7840 10040 8080 10080
rect 6720 10000 7040 10040
rect 7160 10000 7280 10040
rect 7880 10000 8080 10040
rect 6760 9960 7040 10000
rect 7920 9960 8120 10000
rect 6800 9920 7040 9960
rect 7960 9920 8160 9960
rect 6840 9880 7040 9920
rect 8000 9880 8200 9920
rect 6600 9840 6760 9880
rect 6840 9840 7080 9880
rect 6520 9800 6800 9840
rect 6880 9800 7120 9840
rect 8040 9800 8240 9880
rect 6480 9720 6760 9800
rect 6920 9760 7160 9800
rect 8040 9760 8280 9800
rect 6960 9720 7200 9760
rect 8000 9720 8320 9760
rect 6520 9680 6600 9720
rect 7000 9680 7240 9720
rect 7960 9680 8320 9720
rect 7040 9640 7280 9680
rect 7880 9640 8120 9680
rect 8160 9640 8360 9680
rect 7080 9600 7320 9640
rect 7840 9600 8080 9640
rect 6240 9560 6360 9600
rect 7120 9560 7360 9600
rect 7600 9560 8040 9600
rect 8200 9560 8360 9640
rect 6200 8880 6360 9560
rect 7200 9520 7400 9560
rect 7560 9520 8000 9560
rect 7240 9480 7440 9520
rect 7560 9480 7920 9520
rect 7280 9440 7480 9480
rect 7560 9440 7840 9480
rect 6920 9400 7080 9440
rect 7320 9400 7520 9440
rect 6880 9360 7080 9400
rect 7360 9360 7560 9400
rect 6600 9320 7080 9360
rect 6600 9280 7040 9320
rect 7400 9280 7600 9360
rect 6600 9240 6960 9280
rect 7440 9240 7640 9280
rect 6600 9200 6880 9240
rect 7480 9200 7680 9240
rect 7520 9120 7680 9200
rect 7560 9000 7720 9120
rect 8240 9000 8400 9560
rect 7360 8920 7520 8960
rect 7320 8880 7520 8920
rect 5640 8680 5680 8720
rect 5600 8640 5760 8680
rect 6240 8640 6400 8880
rect 7240 8840 7520 8880
rect 7600 8840 7760 9000
rect 8200 8960 8400 9000
rect 8120 8920 8400 8960
rect 8080 8880 8400 8920
rect 8040 8840 8400 8880
rect 6640 8800 6680 8840
rect 7200 8800 7480 8840
rect 6600 8760 6840 8800
rect 7080 8760 7440 8800
rect 6600 8720 7360 8760
rect 6600 8680 7280 8720
rect 6680 8640 7200 8680
rect 5560 8600 5800 8640
rect 5560 8560 5840 8600
rect 5560 8520 5920 8560
rect 6280 8520 6440 8640
rect 7640 8600 7800 8840
rect 7960 8800 8360 8840
rect 7840 8760 8360 8800
rect 7840 8720 8160 8760
rect 7840 8680 8080 8720
rect 7920 8640 7960 8680
rect 7640 8560 7840 8600
rect 5520 8480 6000 8520
rect 5520 8400 5680 8480
rect 5760 8440 6080 8480
rect 6320 8440 6480 8520
rect 5840 8400 6160 8440
rect 6360 8400 6520 8440
rect 5480 8280 5640 8400
rect 5920 8360 6280 8400
rect 5960 8320 6320 8360
rect 6360 8320 6560 8400
rect 6040 8280 6600 8320
rect 5440 8200 5600 8280
rect 6120 8240 6640 8280
rect 6240 8200 6640 8240
rect 6880 8200 7160 8240
rect 7680 8200 7840 8560
rect 5400 8120 5560 8200
rect 6320 8160 7360 8200
rect 5360 8080 5560 8120
rect 6360 8120 7520 8160
rect 6360 8080 7600 8120
rect 5360 8040 5520 8080
rect 6240 8040 6880 8080
rect 7200 8040 7680 8080
rect 7720 8040 7880 8200
rect 5320 8000 5520 8040
rect 6120 8000 6600 8040
rect 7360 8000 7840 8040
rect 5320 7920 5480 8000
rect 6040 7960 6480 8000
rect 7480 7960 7840 8000
rect 5920 7920 6360 7960
rect 7560 7920 7880 7960
rect 5280 7800 5440 7920
rect 5840 7880 6240 7920
rect 7640 7880 7920 7920
rect 5760 7840 6120 7880
rect 7720 7840 7960 7880
rect 8200 7840 8360 8760
rect 5680 7800 6040 7840
rect 7760 7800 8040 7840
rect 5280 7680 5400 7800
rect 5600 7760 5960 7800
rect 7840 7760 8080 7800
rect 5560 7720 5880 7760
rect 7880 7720 8120 7760
rect 5480 7680 5800 7720
rect 7920 7680 8160 7720
rect 8240 7680 8400 7840
rect 5280 7640 5720 7680
rect 7960 7640 8200 7680
rect 8240 7640 8360 7680
rect 5280 7600 5640 7640
rect 8000 7600 8280 7640
rect 5280 7560 5600 7600
rect 8040 7560 8280 7600
rect 5280 7520 5520 7560
rect 8080 7520 8320 7560
rect 5280 7480 5440 7520
rect 8120 7480 8360 7520
rect 5280 7440 5400 7480
rect 8160 7440 8360 7480
rect 5280 7400 5320 7440
rect 6320 7400 6560 7440
rect 8200 7400 8400 7440
rect 6280 7360 6680 7400
rect 6240 7320 6760 7360
rect 8240 7320 8440 7400
rect 6160 7280 6760 7320
rect 8280 7280 8480 7320
rect 6160 7240 6400 7280
rect 6600 7240 6760 7280
rect 8320 7240 8480 7280
rect 6120 7200 6320 7240
rect 6640 7200 6720 7240
rect 8320 7200 8520 7240
rect 6080 7160 6280 7200
rect 8360 7160 8520 7200
rect 6040 7120 6240 7160
rect 8360 7120 8560 7160
rect 6040 7080 6200 7120
rect 6000 7040 6200 7080
rect 7520 7040 7560 7080
rect 8400 7040 8560 7120
rect 6000 6960 6160 7040
rect 7440 6960 7600 7040
rect 8440 6960 8600 7040
rect 5960 6840 6120 6960
rect 7440 6920 7640 6960
rect 8440 6920 8640 6960
rect 7480 6880 7640 6920
rect 7480 6840 7680 6880
rect 8480 6840 8640 6920
rect 5920 6160 6080 6840
rect 7520 6720 7680 6840
rect 8520 6720 8680 6840
rect 7560 6400 7720 6720
rect 8560 6600 8720 6720
rect 8600 6480 8760 6600
rect 7520 6280 7680 6400
rect 8640 6320 8800 6480
rect 7480 6200 7640 6280
rect 7440 6160 7640 6200
rect 8680 6160 8840 6320
rect 3680 5920 3840 5960
rect 3560 5880 3880 5920
rect 3520 5840 3880 5880
rect 3440 5800 3880 5840
rect 5960 5800 6120 6160
rect 7440 6120 7600 6160
rect 7400 6080 7600 6120
rect 7360 6000 7560 6080
rect 7320 5960 7520 6000
rect 8720 5960 8880 6160
rect 7280 5920 7480 5960
rect 7240 5880 7440 5920
rect 7200 5840 7440 5880
rect 7120 5800 7400 5840
rect 3400 5760 3880 5800
rect 3320 5720 3880 5760
rect 3240 5680 3880 5720
rect 3200 5640 3880 5680
rect 3120 5600 3880 5640
rect 3080 5560 3520 5600
rect 3040 5520 3440 5560
rect 3000 5480 3360 5520
rect 1640 5440 1760 5480
rect 3000 5440 3280 5480
rect 1560 4720 1840 5440
rect 3000 5400 3240 5440
rect 3000 5360 3160 5400
rect 3000 5320 3080 5360
rect 920 4680 2480 4720
rect 880 4520 2520 4680
rect 920 4480 2520 4520
rect 960 4440 2480 4480
rect 1560 3760 1840 4440
rect 3600 3800 3880 5600
rect 6000 5240 6120 5800
rect 7080 5760 7360 5800
rect 6960 5720 7280 5760
rect 6880 5680 7240 5720
rect 8760 5680 8920 5960
rect 6760 5640 7200 5680
rect 8800 5640 8920 5680
rect 6640 5600 7080 5640
rect 6560 5560 7000 5600
rect 6480 5520 6920 5560
rect 6440 5480 6760 5520
rect 7120 5480 7400 5520
rect 6400 5440 6680 5480
rect 7040 5440 7480 5480
rect 6360 5400 6600 5440
rect 7000 5400 7560 5440
rect 6280 5360 6560 5400
rect 6920 5360 7600 5400
rect 6240 5320 6480 5360
rect 6880 5320 7640 5360
rect 8800 5320 8960 5640
rect 6200 5280 6440 5320
rect 6840 5280 7680 5320
rect 6160 5240 6400 5280
rect 6800 5240 7320 5280
rect 7520 5240 7720 5280
rect 6000 5200 6360 5240
rect 5960 5160 6320 5200
rect 6760 5160 7240 5240
rect 7560 5200 7760 5240
rect 7600 5160 7760 5200
rect 5960 5120 6280 5160
rect 5960 5080 6240 5120
rect 6720 5080 7200 5160
rect 7640 5120 7800 5160
rect 5960 5040 6200 5080
rect 6680 5040 7200 5080
rect 7680 5080 7800 5120
rect 7680 5040 7840 5080
rect 5920 5000 6200 5040
rect 5920 4960 6160 5000
rect 5920 4880 6120 4960
rect 6640 4920 7200 5040
rect 7720 4960 7840 5040
rect 8840 4960 9000 5320
rect 5880 4800 6080 4880
rect 6600 4840 7240 4920
rect 7720 4880 7880 4960
rect 7680 4840 7880 4880
rect 6600 4800 7280 4840
rect 7640 4800 7880 4840
rect 5880 4720 6040 4800
rect 6600 4760 7440 4800
rect 7520 4760 7880 4800
rect 5920 4680 6000 4720
rect 6560 4600 7880 4760
rect 8880 4920 9000 4960
rect 11080 5000 11200 5040
rect 11080 4960 11320 5000
rect 11080 4920 11400 4960
rect 8880 4680 9040 4920
rect 11080 4880 11440 4920
rect 11200 4840 11480 4880
rect 11280 4800 11520 4840
rect 11360 4760 11560 4800
rect 11400 4720 11560 4760
rect 8880 4640 9080 4680
rect 6600 4400 7880 4600
rect 8920 4600 9080 4640
rect 8920 4560 9120 4600
rect 10920 4560 11040 4600
rect 8960 4520 9120 4560
rect 10880 4520 11080 4560
rect 8960 4480 9160 4520
rect 6640 4360 7880 4400
rect 6640 4320 7840 4360
rect 6680 4240 7840 4320
rect 9000 4240 9160 4480
rect 10880 4400 11040 4520
rect 11440 4480 11600 4720
rect 11440 4440 11640 4480
rect 11480 4400 11640 4440
rect 10840 4360 11040 4400
rect 10800 4320 11040 4360
rect 11520 4320 11680 4400
rect 10760 4280 11000 4320
rect 10720 4240 10920 4280
rect 6720 4200 7840 4240
rect 9040 4200 9160 4240
rect 10680 4200 10880 4240
rect 6760 4120 7800 4200
rect 6800 4080 7760 4120
rect 6840 4040 7760 4080
rect 6880 4000 7720 4040
rect 6920 3960 7680 4000
rect 7000 3920 7640 3960
rect 9040 3920 9200 4200
rect 10640 4160 10840 4200
rect 10640 4120 10800 4160
rect 10600 4040 10760 4120
rect 11560 4080 11720 4320
rect 11520 4040 11720 4080
rect 10600 4000 10720 4040
rect 11480 4000 11680 4040
rect 7040 3880 7560 3920
rect 7120 3840 7480 3880
rect 3560 3760 3880 3800
rect 1600 3720 1800 3760
rect 3040 3720 4360 3760
rect 3000 3560 4400 3720
rect 9080 3680 9240 3920
rect 10560 3760 10720 4000
rect 11440 3960 11640 4000
rect 11360 3920 11640 3960
rect 11320 3880 11560 3920
rect 11240 3840 11520 3880
rect 11240 3800 11480 3840
rect 11240 3760 11440 3800
rect 10600 3680 10760 3760
rect 11280 3720 11480 3760
rect 11320 3680 11520 3720
rect 3040 3520 4360 3560
rect 9120 3480 9280 3680
rect 10600 3640 10800 3680
rect 11360 3640 11520 3680
rect 10640 3560 10840 3640
rect 11400 3560 11560 3640
rect 10600 3480 10840 3560
rect 5920 3360 6040 3400
rect 9160 3360 9320 3480
rect 10560 3440 10760 3480
rect 10560 3400 10720 3440
rect 10520 3360 10720 3400
rect 5880 3280 6040 3360
rect 5840 3240 6040 3280
rect 9200 3280 9360 3360
rect 9200 3240 9400 3280
rect 10520 3240 10680 3360
rect 11440 3320 11600 3560
rect 11400 3280 11600 3320
rect 11400 3240 11560 3280
rect 5800 3200 6000 3240
rect 9240 3200 9400 3240
rect 5800 3160 5960 3200
rect 9240 3160 9440 3200
rect 10480 3160 10640 3240
rect 11360 3200 11560 3240
rect 11280 3160 11520 3200
rect 5760 3120 5960 3160
rect 9280 3120 9440 3160
rect 5760 3080 5920 3120
rect 9280 3080 9480 3120
rect 5720 3040 5920 3080
rect 9320 3040 9480 3080
rect 5720 3000 5880 3040
rect 9320 3000 9520 3040
rect 10520 3000 10680 3160
rect 11240 3120 11480 3160
rect 11200 3080 11440 3120
rect 11240 3040 11400 3080
rect 11240 3000 11360 3040
rect 5680 2960 5880 3000
rect 9360 2960 9520 3000
rect 10560 2960 10720 3000
rect 5680 2840 5840 2960
rect 9360 2920 9560 2960
rect 10560 2920 10760 2960
rect 9400 2880 9640 2920
rect 10600 2880 10800 2920
rect 9440 2840 9760 2880
rect 10600 2840 10840 2880
rect 5640 2720 5800 2840
rect 9480 2800 9880 2840
rect 10640 2800 10920 2840
rect 9520 2760 10040 2800
rect 10680 2760 10960 2800
rect 9600 2720 10160 2760
rect 10720 2720 11000 2760
rect 5680 2680 5800 2720
rect 9720 2680 10280 2720
rect 10800 2680 10960 2720
rect 5680 2560 5840 2680
rect 9840 2640 10320 2680
rect 10880 2640 10920 2680
rect 10000 2600 10400 2640
rect 10160 2560 10440 2600
rect 5720 2520 5880 2560
rect 10240 2520 10520 2560
rect 5720 2480 5920 2520
rect 10320 2480 10560 2520
rect 5760 2440 5920 2480
rect 10360 2440 10600 2480
rect 5720 2400 5960 2440
rect 10440 2400 10640 2440
rect 5680 2360 6000 2400
rect 10480 2360 10680 2400
rect 5600 2320 6040 2360
rect 10520 2320 10720 2360
rect 5560 2280 6120 2320
rect 10560 2280 10720 2320
rect 5480 2240 5760 2280
rect 5920 2240 6160 2280
rect 7320 2240 7360 2280
rect 10560 2240 10760 2280
rect 5440 2200 5720 2240
rect 5960 2200 6240 2240
rect 7240 2200 7400 2240
rect 10600 2200 10760 2240
rect 5400 2160 5640 2200
rect 6000 2160 6360 2200
rect 7200 2160 7400 2200
rect 5320 2120 5600 2160
rect 6080 2120 6440 2160
rect 7160 2120 7400 2160
rect 10200 2120 10280 2160
rect 10640 2120 10800 2200
rect 5280 2080 5560 2120
rect 6160 2080 6600 2120
rect 7080 2080 7360 2120
rect 5280 2040 5480 2080
rect 6240 2040 7320 2080
rect 5280 2000 5440 2040
rect 6320 2000 7240 2040
rect 5280 1960 5400 2000
rect 6440 1960 7160 2000
rect 5280 1920 5360 1960
rect 6600 1920 7040 1960
rect 10160 1920 10320 2120
rect 10680 1960 10840 2120
rect 5280 1880 5320 1920
rect 6840 1880 7040 1920
rect 6880 1840 7080 1880
rect 10120 1840 10280 1920
rect 10720 1880 10840 1960
rect 6880 1800 7120 1840
rect 10080 1800 10280 1840
rect 6920 1760 7160 1800
rect 10080 1760 10240 1800
rect 6960 1720 7200 1760
rect 10080 1720 10200 1760
rect 7000 1680 7240 1720
rect 8800 1680 8920 1720
rect 10120 1680 10160 1720
rect 7040 1640 7320 1680
rect 8800 1640 8960 1680
rect 10680 1640 10840 1880
rect 7080 1600 7360 1640
rect 8800 1600 9040 1640
rect 7160 1560 7400 1600
rect 8840 1560 9080 1600
rect 10640 1560 10800 1640
rect 7200 1520 7480 1560
rect 8880 1520 9120 1560
rect 10600 1520 10800 1560
rect 7240 1480 7520 1520
rect 8920 1480 9160 1520
rect 7320 1440 7600 1480
rect 8960 1440 9240 1480
rect 10600 1440 10760 1520
rect 7360 1400 7680 1440
rect 9040 1400 9280 1440
rect 7440 1360 7720 1400
rect 9080 1360 9320 1400
rect 10560 1360 10720 1440
rect 7480 1320 7800 1360
rect 9120 1320 9360 1360
rect 10520 1320 10720 1360
rect 7560 1280 7880 1320
rect 9160 1280 9400 1320
rect 10480 1280 10680 1320
rect 7640 1240 7960 1280
rect 9240 1240 9440 1280
rect 10480 1240 10640 1280
rect 7680 1200 8040 1240
rect 9280 1200 9520 1240
rect 10440 1200 10640 1240
rect 7760 1160 8120 1200
rect 9320 1160 9560 1200
rect 10400 1160 10600 1200
rect 7840 1120 8200 1160
rect 9360 1120 9600 1160
rect 10360 1120 10560 1160
rect 7920 1080 8320 1120
rect 9400 1080 9640 1120
rect 10320 1080 10520 1120
rect 8000 1040 8400 1080
rect 9440 1040 9720 1080
rect 10280 1040 10520 1080
rect 8080 1000 8520 1040
rect 9400 1000 9760 1040
rect 10240 1000 10480 1040
rect 8160 960 8640 1000
rect 9320 960 9840 1000
rect 10200 960 10440 1000
rect 8280 920 8920 960
rect 9120 920 9560 960
rect 9640 920 9880 960
rect 10160 920 10400 960
rect 8360 880 9480 920
rect 9680 880 9960 920
rect 10120 880 10360 920
rect 8480 840 9440 880
rect 9720 840 10320 880
rect 8640 800 9360 840
rect 9800 800 10280 840
rect 8920 760 9160 800
rect 9880 760 10240 800
rect 9920 720 10160 760
<< end >>
