magic
tech sky130A
magscale 1 2
timestamp 1754836895
<< locali >>
rect 10800 9100 13200 10600
rect 12500 8000 13200 9100
rect 10700 6500 13200 8000
rect 14300 9100 16900 10900
rect 23800 10800 25800 10900
rect 14300 8000 15100 9100
rect 14300 6500 16800 8000
rect 23800 7500 23900 10800
rect 25600 7500 25800 10800
rect 23800 7200 25800 7500
rect 23800 6200 23900 7200
rect 22900 3900 23900 6200
rect 25600 3900 25800 7200
rect 22900 3600 25800 3900
rect 12264 2904 15316 3096
rect 12500 600 15100 2904
rect 12500 100 14200 600
rect 15238 170 15650 230
rect 22900 226 23900 3600
rect 25600 232 25800 3600
rect 24877 226 25800 232
rect 14384 70 14796 76
rect 14384 -110 14390 70
rect 14570 -110 14796 70
rect 16360 -70 16462 -10
rect 16632 -108 17028 68
rect 14384 -116 14796 -110
rect 16852 -218 17028 -108
rect 16852 -382 16858 -218
rect 17022 -382 17028 -218
rect 16852 -388 17028 -382
rect 22900 -14 25800 226
rect 22900 -240 23900 -14
rect 22900 -480 24404 -240
rect 14000 -4580 14600 -600
rect 15618 -730 15630 -670
rect 15570 -850 15630 -730
rect 22900 -800 23900 -480
rect 17400 -980 23900 -800
rect 17400 -1220 22580 -980
rect 22808 -1220 23900 -980
rect 16170 -3382 16230 -3270
rect 17400 -3300 23900 -1220
rect 25600 -3300 25800 -14
rect 17400 -3500 25800 -3300
rect 14770 -4130 14880 -4070
rect 17400 -4200 23000 -3500
rect 13940 -4600 14600 -4580
rect 13800 -4700 14600 -4600
rect 15930 -4656 15990 -4490
rect 13800 -5012 14180 -4700
rect 15930 -4704 15936 -4656
rect 15984 -4704 15990 -4656
rect 15930 -4710 15990 -4704
rect 17400 -4900 19100 -4200
rect 13800 -5584 14000 -5012
rect 15100 -5504 19100 -4900
rect 13800 -5924 14180 -5584
rect 15012 -5780 19100 -5504
rect 13800 -6420 14000 -5924
rect 15012 -5936 15348 -5780
rect 15082 -5944 15348 -5936
rect 15512 -5944 19100 -5780
rect 15082 -5950 19100 -5944
rect 15100 -6404 19100 -5950
rect 13800 -6604 14180 -6420
rect 15012 -6604 19100 -6404
rect 13800 -6610 19100 -6604
rect 13800 -6790 14378 -6610
rect 14558 -6790 19100 -6610
rect 13800 -7100 19100 -6790
<< viali >>
rect 24164 10320 24404 10560
rect 25076 10320 25316 10560
rect 24164 6720 24404 6960
rect 25076 6720 25316 6960
rect 15190 170 15238 230
rect 24164 3120 24392 3360
rect 25088 3120 25316 3360
rect 14390 -110 14570 70
rect 16462 -70 16510 -10
rect 16858 -382 17022 -218
rect 25088 -480 25316 -240
rect 15570 -730 15618 -670
rect 22580 -1220 22808 -980
rect 16170 -3430 16230 -3382
rect 15936 -4704 15984 -4656
rect 15348 -5944 15512 -5780
rect 14378 -6790 14558 -6610
<< metal1 >>
rect 4500 10920 23700 11000
rect 4500 10600 23720 10920
rect 13850 9204 13856 9396
rect 14048 9204 14054 9396
rect 14300 456 14700 10600
rect 23480 10560 23720 10600
rect 24140 10560 24420 10580
rect 23480 10320 24164 10560
rect 24404 10320 24420 10560
rect 24140 10300 24420 10320
rect 25060 10560 25520 10580
rect 25060 10320 25076 10560
rect 25316 10320 25520 10560
rect 25060 10300 25520 10320
rect 25280 6980 25520 10300
rect 23980 6960 24420 6980
rect 23980 6720 24164 6960
rect 24404 6720 24420 6960
rect 23980 6700 24420 6720
rect 25060 6960 25520 6980
rect 25060 6720 25076 6960
rect 25316 6720 25520 6960
rect 25060 6700 25520 6720
rect 23980 3372 24220 6700
rect 25316 3762 25520 3768
rect 25316 3372 25520 3558
rect 23980 3360 24398 3372
rect 14850 3150 15470 3210
rect 14850 590 14910 3150
rect 23980 3120 24164 3360
rect 24392 3120 24398 3360
rect 24158 3108 24398 3120
rect 25082 3360 25520 3372
rect 25082 3120 25088 3360
rect 25316 3120 25520 3360
rect 25082 3108 25520 3120
rect 14850 530 16516 590
rect 14300 264 14964 456
rect 15156 264 15162 456
rect 14300 70 14700 264
rect 14300 -110 14390 70
rect 14570 -110 14700 70
rect 14300 -200 14700 -110
rect 15184 230 15244 242
rect 15184 170 15190 230
rect 15238 170 15244 230
rect 15184 -210 15244 170
rect 16456 -10 16516 530
rect 16456 -70 16462 -10
rect 16510 -70 16516 -10
rect 16456 -82 16516 -70
rect 15184 -276 15244 -270
rect 16212 -212 16388 -206
rect 16388 -218 17034 -212
rect 16388 -382 16858 -218
rect 17022 -382 17034 -218
rect 25280 -228 25520 3108
rect 16388 -388 17034 -382
rect 25082 -240 25520 -228
rect 16212 -394 16388 -388
rect 25082 -480 25088 -240
rect 25316 -480 25520 -240
rect 25082 -492 25322 -480
rect 15564 -670 15624 -658
rect 15064 -730 15070 -670
rect 15130 -730 15570 -670
rect 15618 -730 15624 -670
rect 15564 -742 15624 -730
rect 22574 -980 22814 -968
rect 22174 -1220 22180 -980
rect 22420 -1220 22580 -980
rect 22808 -1220 22814 -980
rect 22574 -1232 22814 -1220
rect 16158 -3382 16242 -3376
rect 16158 -3430 16170 -3382
rect 16230 -3430 16242 -3382
rect 16158 -3436 16242 -3430
rect 16170 -3470 16230 -3436
rect 16170 -3536 16230 -3530
rect 14700 -4650 14760 -3910
rect 14700 -4656 15996 -4650
rect 14700 -4704 15936 -4656
rect 15984 -4704 15996 -4656
rect 14700 -4710 15996 -4704
rect 14230 -4852 14320 -4840
rect 14230 -4916 14244 -4852
rect 14308 -4916 14320 -4852
rect 14230 -4930 14320 -4916
rect 14628 -5044 15284 -4852
rect 15476 -5044 15482 -4852
rect 14244 -5892 14308 -5508
rect 14372 -5936 14564 -5148
rect 14628 -5936 14820 -5244
rect 15336 -5650 15342 -5474
rect 15518 -5650 15524 -5474
rect 15342 -5780 15518 -5650
rect 15342 -5944 15348 -5780
rect 15512 -5944 15518 -5780
rect 15342 -5956 15518 -5944
rect 14372 -6610 14564 -6104
rect 14372 -6790 14378 -6610
rect 14558 -6790 14564 -6610
rect 14372 -6802 14564 -6790
<< via1 >>
rect 13856 9204 14048 9396
rect 25316 3558 25520 3762
rect 14964 264 15156 456
rect 15184 -270 15244 -210
rect 16212 -388 16388 -212
rect 15070 -730 15130 -670
rect 22180 -1220 22420 -980
rect 16170 -3530 16230 -3470
rect 14244 -4916 14308 -4852
rect 15284 -5044 15476 -4852
rect 15342 -5650 15518 -5474
<< metal2 >>
rect 13856 9396 14048 9402
rect 14048 9204 14634 9396
rect 14816 9204 14825 9396
rect 13856 9198 14048 9204
rect 14720 6442 23620 6580
rect 14720 6340 23622 6442
rect 14720 5700 14960 6340
rect 23380 3762 23622 6340
rect 23380 3560 25316 3762
rect 23418 3558 25316 3560
rect 25520 3558 25526 3762
rect 9230 1420 14630 1480
rect 14964 456 15156 462
rect 15156 264 15334 456
rect 15516 264 15525 456
rect 14964 258 15156 264
rect 15178 -270 15184 -210
rect 15244 -270 15250 -210
rect 15884 -217 16212 -212
rect 15184 -570 15244 -270
rect 15880 -383 15889 -217
rect 16055 -383 16212 -217
rect 15884 -388 16212 -383
rect 16388 -388 16394 -212
rect 15184 -630 16430 -570
rect 15070 -670 15130 -664
rect 14270 -692 15070 -670
rect 14244 -730 15070 -692
rect 14244 -4840 14308 -730
rect 15070 -736 15130 -730
rect 16370 -3470 16430 -630
rect 22180 -980 22420 -974
rect 21771 -1220 21780 -980
rect 22010 -1220 22180 -980
rect 22180 -1226 22420 -1220
rect 16164 -3530 16170 -3470
rect 16230 -3530 16430 -3470
rect 14230 -4852 14320 -4840
rect 14230 -4916 14244 -4852
rect 14308 -4916 14320 -4852
rect 14230 -4930 14320 -4916
rect 15284 -4852 15476 -4846
rect 15476 -5044 15874 -4852
rect 16056 -5044 16065 -4852
rect 15284 -5050 15476 -5044
rect 15342 -5115 15518 -5110
rect 15338 -5281 15347 -5115
rect 15513 -5281 15522 -5115
rect 15342 -5474 15518 -5281
rect 15342 -5656 15518 -5650
<< via2 >>
rect 14634 9204 14816 9396
rect 15334 264 15516 456
rect 15889 -383 16055 -217
rect 21780 -1220 22010 -980
rect 15874 -5044 16056 -4852
rect 15347 -5281 15513 -5115
<< metal3 >>
rect 14629 9396 14821 9401
rect 14629 9204 14634 9396
rect 14816 9204 14821 9396
rect 14629 6316 14821 9204
rect 14629 6124 18536 6316
rect 15329 456 15521 461
rect 15329 264 15334 456
rect 15516 264 15521 456
rect 15329 -424 15521 264
rect 15884 -217 16060 -24
rect 15884 -383 15889 -217
rect 16055 -383 16060 -217
rect 15884 -388 16060 -383
rect 15329 -512 15836 -424
rect 15329 -616 15896 -512
rect 15720 -1588 15896 -616
rect 18344 -1496 18536 6124
rect 21775 -980 22015 -975
rect 21374 -1220 21380 -980
rect 21618 -1220 21780 -980
rect 22010 -1220 22015 -980
rect 21775 -1225 22015 -1220
rect 16904 -3596 18096 -3404
rect 15180 -5110 15356 -4344
rect 15869 -4852 16061 -4847
rect 16904 -4852 17096 -3596
rect 15869 -5044 15874 -4852
rect 16056 -5044 17096 -4852
rect 15869 -5049 16061 -5044
rect 15180 -5115 15518 -5110
rect 15180 -5281 15347 -5115
rect 15513 -5281 15518 -5115
rect 15180 -5286 15518 -5281
<< via3 >>
rect 21380 -1220 21618 -980
<< metal4 >>
rect 21379 -980 21619 -979
rect 21379 -1220 21380 -980
rect 21618 -1220 21619 -980
rect 21379 -1380 21619 -1220
rect 20080 -1620 21619 -1380
use JNWATR_NCH_2C1F2 JNWATR_NCH_2C1F2_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 14084 0 1 -6572
box -184 -128 1208 928
use JNWATR_NCH_2C1F2 JNWATR_NCH_2C1F2_1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 14084 0 1 -5612
box -184 -128 1208 928
use JNWTR_BFX1_CV x3 ../JNW_TR_SKY130A
timestamp 1754771195
transform -1 0 16690 0 1 -200
box -150 -120 2130 600
use amplifier_rev2 x4 ../JNW_GR07_SKY130A
timestamp 1754836895
transform -1 0 22000 0 1 2600
box -1600 -3400 7200 8300
use JNWTR_DFRNQNX1_CV x5 ../JNW_TR_SKY130A
timestamp 1754771195
transform 1 0 14550 0 1 -4580
box -150 -120 2130 3960
use JNWTR_RPPO4 x6 ../JNW_TR_SKY130A
timestamp 1754770625
transform -1 0 25680 0 1 7400
box 0 0 1880 3440
use JNWTR_CAPX4 x7 ../JNW_TR_SKY130A
timestamp 1754836895
transform 1 0 17320 0 1 -3800
box 480 0 3120 2640
use JNWTR_RPPO4 x8 ../JNW_TR_SKY130A
timestamp 1754770625
transform 1 0 23800 0 1 -3400
box 0 0 1880 3440
use JNWTR_RPPO4 x9 ../JNW_TR_SKY130A
timestamp 1754770625
transform -1 0 25680 0 1 200
box 0 0 1880 3440
use JNWTR_RPPO4 x10 ../JNW_TR_SKY130A
timestamp 1754770625
transform 1 0 23800 0 1 3800
box 0 0 1880 3440
use temp_to_current_rev2 x11 ../JNW_GR07_SKY130A
timestamp 1754836895
transform 1 0 4600 0 1 2800
box -600 -10800 9920 8100
<< labels >>
flabel space 9000 -8000 9500 -7500 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel metal1 14924 10684 15116 10876 0 FreeSans 1600 0 0 0 VDD
port 13 nsew
flabel metal2 14270 -4852 14308 -670 0 FreeSans 1600 0 0 0 PWM
port 15 nsew
flabel locali 14770 -4130 14880 -4070 0 FreeSans 1600 0 0 0 CLK
port 16 nsew
flabel locali 15012 -6796 15204 -6604 0 FreeSans 1600 0 0 0 VSS
port 17 nsew
<< properties >>
string FIXED_BBOX 3950 -8076 25750 10920
<< end >>
