magic
tech sky130A
magscale 1 2
timestamp 1757256469
<< nwell >>
rect -1809 -362 1809 362
<< mvpmos >>
rect -1551 -64 -1451 136
rect -1393 -64 -1293 136
rect -1235 -64 -1135 136
rect -1077 -64 -977 136
rect -919 -64 -819 136
rect -761 -64 -661 136
rect -603 -64 -503 136
rect -445 -64 -345 136
rect -287 -64 -187 136
rect -129 -64 -29 136
rect 29 -64 129 136
rect 187 -64 287 136
rect 345 -64 445 136
rect 503 -64 603 136
rect 661 -64 761 136
rect 819 -64 919 136
rect 977 -64 1077 136
rect 1135 -64 1235 136
rect 1293 -64 1393 136
rect 1451 -64 1551 136
<< mvpdiff >>
rect -1609 124 -1551 136
rect -1609 -52 -1597 124
rect -1563 -52 -1551 124
rect -1609 -64 -1551 -52
rect -1451 124 -1393 136
rect -1451 -52 -1439 124
rect -1405 -52 -1393 124
rect -1451 -64 -1393 -52
rect -1293 124 -1235 136
rect -1293 -52 -1281 124
rect -1247 -52 -1235 124
rect -1293 -64 -1235 -52
rect -1135 124 -1077 136
rect -1135 -52 -1123 124
rect -1089 -52 -1077 124
rect -1135 -64 -1077 -52
rect -977 124 -919 136
rect -977 -52 -965 124
rect -931 -52 -919 124
rect -977 -64 -919 -52
rect -819 124 -761 136
rect -819 -52 -807 124
rect -773 -52 -761 124
rect -819 -64 -761 -52
rect -661 124 -603 136
rect -661 -52 -649 124
rect -615 -52 -603 124
rect -661 -64 -603 -52
rect -503 124 -445 136
rect -503 -52 -491 124
rect -457 -52 -445 124
rect -503 -64 -445 -52
rect -345 124 -287 136
rect -345 -52 -333 124
rect -299 -52 -287 124
rect -345 -64 -287 -52
rect -187 124 -129 136
rect -187 -52 -175 124
rect -141 -52 -129 124
rect -187 -64 -129 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 129 124 187 136
rect 129 -52 141 124
rect 175 -52 187 124
rect 129 -64 187 -52
rect 287 124 345 136
rect 287 -52 299 124
rect 333 -52 345 124
rect 287 -64 345 -52
rect 445 124 503 136
rect 445 -52 457 124
rect 491 -52 503 124
rect 445 -64 503 -52
rect 603 124 661 136
rect 603 -52 615 124
rect 649 -52 661 124
rect 603 -64 661 -52
rect 761 124 819 136
rect 761 -52 773 124
rect 807 -52 819 124
rect 761 -64 819 -52
rect 919 124 977 136
rect 919 -52 931 124
rect 965 -52 977 124
rect 919 -64 977 -52
rect 1077 124 1135 136
rect 1077 -52 1089 124
rect 1123 -52 1135 124
rect 1077 -64 1135 -52
rect 1235 124 1293 136
rect 1235 -52 1247 124
rect 1281 -52 1293 124
rect 1235 -64 1293 -52
rect 1393 124 1451 136
rect 1393 -52 1405 124
rect 1439 -52 1451 124
rect 1393 -64 1451 -52
rect 1551 124 1609 136
rect 1551 -52 1563 124
rect 1597 -52 1609 124
rect 1551 -64 1609 -52
<< mvpdiffc >>
rect -1597 -52 -1563 124
rect -1439 -52 -1405 124
rect -1281 -52 -1247 124
rect -1123 -52 -1089 124
rect -965 -52 -931 124
rect -807 -52 -773 124
rect -649 -52 -615 124
rect -491 -52 -457 124
rect -333 -52 -299 124
rect -175 -52 -141 124
rect -17 -52 17 124
rect 141 -52 175 124
rect 299 -52 333 124
rect 457 -52 491 124
rect 615 -52 649 124
rect 773 -52 807 124
rect 931 -52 965 124
rect 1089 -52 1123 124
rect 1247 -52 1281 124
rect 1405 -52 1439 124
rect 1563 -52 1597 124
<< mvnsubdiff >>
rect -1743 284 1743 296
rect -1743 250 -1635 284
rect 1635 250 1743 284
rect -1743 238 1743 250
rect -1743 188 -1685 238
rect -1743 -188 -1731 188
rect -1697 -188 -1685 188
rect 1685 188 1743 238
rect -1743 -238 -1685 -188
rect 1685 -188 1697 188
rect 1731 -188 1743 188
rect 1685 -238 1743 -188
rect -1743 -250 1743 -238
rect -1743 -284 -1635 -250
rect 1635 -284 1743 -250
rect -1743 -296 1743 -284
<< mvnsubdiffcont >>
rect -1635 250 1635 284
rect -1731 -188 -1697 188
rect 1697 -188 1731 188
rect -1635 -284 1635 -250
<< poly >>
rect -1551 136 -1451 162
rect -1393 136 -1293 162
rect -1235 136 -1135 162
rect -1077 136 -977 162
rect -919 136 -819 162
rect -761 136 -661 162
rect -603 136 -503 162
rect -445 136 -345 162
rect -287 136 -187 162
rect -129 136 -29 162
rect 29 136 129 162
rect 187 136 287 162
rect 345 136 445 162
rect 503 136 603 162
rect 661 136 761 162
rect 819 136 919 162
rect 977 136 1077 162
rect 1135 136 1235 162
rect 1293 136 1393 162
rect 1451 136 1551 162
rect -1551 -111 -1451 -64
rect -1551 -145 -1535 -111
rect -1467 -145 -1451 -111
rect -1551 -161 -1451 -145
rect -1393 -111 -1293 -64
rect -1393 -145 -1377 -111
rect -1309 -145 -1293 -111
rect -1393 -161 -1293 -145
rect -1235 -111 -1135 -64
rect -1235 -145 -1219 -111
rect -1151 -145 -1135 -111
rect -1235 -161 -1135 -145
rect -1077 -111 -977 -64
rect -1077 -145 -1061 -111
rect -993 -145 -977 -111
rect -1077 -161 -977 -145
rect -919 -111 -819 -64
rect -919 -145 -903 -111
rect -835 -145 -819 -111
rect -919 -161 -819 -145
rect -761 -111 -661 -64
rect -761 -145 -745 -111
rect -677 -145 -661 -111
rect -761 -161 -661 -145
rect -603 -111 -503 -64
rect -603 -145 -587 -111
rect -519 -145 -503 -111
rect -603 -161 -503 -145
rect -445 -111 -345 -64
rect -445 -145 -429 -111
rect -361 -145 -345 -111
rect -445 -161 -345 -145
rect -287 -111 -187 -64
rect -287 -145 -271 -111
rect -203 -145 -187 -111
rect -287 -161 -187 -145
rect -129 -111 -29 -64
rect -129 -145 -113 -111
rect -45 -145 -29 -111
rect -129 -161 -29 -145
rect 29 -111 129 -64
rect 29 -145 45 -111
rect 113 -145 129 -111
rect 29 -161 129 -145
rect 187 -111 287 -64
rect 187 -145 203 -111
rect 271 -145 287 -111
rect 187 -161 287 -145
rect 345 -111 445 -64
rect 345 -145 361 -111
rect 429 -145 445 -111
rect 345 -161 445 -145
rect 503 -111 603 -64
rect 503 -145 519 -111
rect 587 -145 603 -111
rect 503 -161 603 -145
rect 661 -111 761 -64
rect 661 -145 677 -111
rect 745 -145 761 -111
rect 661 -161 761 -145
rect 819 -111 919 -64
rect 819 -145 835 -111
rect 903 -145 919 -111
rect 819 -161 919 -145
rect 977 -111 1077 -64
rect 977 -145 993 -111
rect 1061 -145 1077 -111
rect 977 -161 1077 -145
rect 1135 -111 1235 -64
rect 1135 -145 1151 -111
rect 1219 -145 1235 -111
rect 1135 -161 1235 -145
rect 1293 -111 1393 -64
rect 1293 -145 1309 -111
rect 1377 -145 1393 -111
rect 1293 -161 1393 -145
rect 1451 -111 1551 -64
rect 1451 -145 1467 -111
rect 1535 -145 1551 -111
rect 1451 -161 1551 -145
<< polycont >>
rect -1535 -145 -1467 -111
rect -1377 -145 -1309 -111
rect -1219 -145 -1151 -111
rect -1061 -145 -993 -111
rect -903 -145 -835 -111
rect -745 -145 -677 -111
rect -587 -145 -519 -111
rect -429 -145 -361 -111
rect -271 -145 -203 -111
rect -113 -145 -45 -111
rect 45 -145 113 -111
rect 203 -145 271 -111
rect 361 -145 429 -111
rect 519 -145 587 -111
rect 677 -145 745 -111
rect 835 -145 903 -111
rect 993 -145 1061 -111
rect 1151 -145 1219 -111
rect 1309 -145 1377 -111
rect 1467 -145 1535 -111
<< locali >>
rect -1731 250 -1635 284
rect 1635 250 1731 284
rect -1731 188 -1697 250
rect 1697 188 1731 250
rect -1597 124 -1563 140
rect -1597 -68 -1563 -52
rect -1439 124 -1405 140
rect -1439 -68 -1405 -52
rect -1281 124 -1247 140
rect -1281 -68 -1247 -52
rect -1123 124 -1089 140
rect -1123 -68 -1089 -52
rect -965 124 -931 140
rect -965 -68 -931 -52
rect -807 124 -773 140
rect -807 -68 -773 -52
rect -649 124 -615 140
rect -649 -68 -615 -52
rect -491 124 -457 140
rect -491 -68 -457 -52
rect -333 124 -299 140
rect -333 -68 -299 -52
rect -175 124 -141 140
rect -175 -68 -141 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 141 124 175 140
rect 141 -68 175 -52
rect 299 124 333 140
rect 299 -68 333 -52
rect 457 124 491 140
rect 457 -68 491 -52
rect 615 124 649 140
rect 615 -68 649 -52
rect 773 124 807 140
rect 773 -68 807 -52
rect 931 124 965 140
rect 931 -68 965 -52
rect 1089 124 1123 140
rect 1089 -68 1123 -52
rect 1247 124 1281 140
rect 1247 -68 1281 -52
rect 1405 124 1439 140
rect 1405 -68 1439 -52
rect 1563 124 1597 140
rect 1563 -68 1597 -52
rect -1551 -145 -1535 -111
rect -1467 -145 -1451 -111
rect -1393 -145 -1377 -111
rect -1309 -145 -1293 -111
rect -1235 -145 -1219 -111
rect -1151 -145 -1135 -111
rect -1077 -145 -1061 -111
rect -993 -145 -977 -111
rect -919 -145 -903 -111
rect -835 -145 -819 -111
rect -761 -145 -745 -111
rect -677 -145 -661 -111
rect -603 -145 -587 -111
rect -519 -145 -503 -111
rect -445 -145 -429 -111
rect -361 -145 -345 -111
rect -287 -145 -271 -111
rect -203 -145 -187 -111
rect -129 -145 -113 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 113 -145 129 -111
rect 187 -145 203 -111
rect 271 -145 287 -111
rect 345 -145 361 -111
rect 429 -145 445 -111
rect 503 -145 519 -111
rect 587 -145 603 -111
rect 661 -145 677 -111
rect 745 -145 761 -111
rect 819 -145 835 -111
rect 903 -145 919 -111
rect 977 -145 993 -111
rect 1061 -145 1077 -111
rect 1135 -145 1151 -111
rect 1219 -145 1235 -111
rect 1293 -145 1309 -111
rect 1377 -145 1393 -111
rect 1451 -145 1467 -111
rect 1535 -145 1551 -111
rect -1731 -250 -1697 -188
rect 1697 -250 1731 -188
rect -1731 -284 -1635 -250
rect 1635 -284 1731 -250
<< viali >>
rect -1597 -52 -1563 124
rect -1439 -52 -1405 124
rect -1281 -52 -1247 124
rect -1123 -52 -1089 124
rect -965 -52 -931 124
rect -807 -52 -773 124
rect -649 -52 -615 124
rect -491 -52 -457 124
rect -333 -52 -299 124
rect -175 -52 -141 124
rect -17 -52 17 124
rect 141 -52 175 124
rect 299 -52 333 124
rect 457 -52 491 124
rect 615 -52 649 124
rect 773 -52 807 124
rect 931 -52 965 124
rect 1089 -52 1123 124
rect 1247 -52 1281 124
rect 1405 -52 1439 124
rect 1563 -52 1597 124
rect -1535 -145 -1467 -111
rect -1377 -145 -1309 -111
rect -1219 -145 -1151 -111
rect -1061 -145 -993 -111
rect -903 -145 -835 -111
rect -745 -145 -677 -111
rect -587 -145 -519 -111
rect -429 -145 -361 -111
rect -271 -145 -203 -111
rect -113 -145 -45 -111
rect 45 -145 113 -111
rect 203 -145 271 -111
rect 361 -145 429 -111
rect 519 -145 587 -111
rect 677 -145 745 -111
rect 835 -145 903 -111
rect 993 -145 1061 -111
rect 1151 -145 1219 -111
rect 1309 -145 1377 -111
rect 1467 -145 1535 -111
<< metal1 >>
rect -1603 124 -1557 136
rect -1603 -52 -1597 124
rect -1563 -52 -1557 124
rect -1603 -64 -1557 -52
rect -1445 124 -1399 136
rect -1445 -52 -1439 124
rect -1405 -52 -1399 124
rect -1445 -64 -1399 -52
rect -1287 124 -1241 136
rect -1287 -52 -1281 124
rect -1247 -52 -1241 124
rect -1287 -64 -1241 -52
rect -1129 124 -1083 136
rect -1129 -52 -1123 124
rect -1089 -52 -1083 124
rect -1129 -64 -1083 -52
rect -971 124 -925 136
rect -971 -52 -965 124
rect -931 -52 -925 124
rect -971 -64 -925 -52
rect -813 124 -767 136
rect -813 -52 -807 124
rect -773 -52 -767 124
rect -813 -64 -767 -52
rect -655 124 -609 136
rect -655 -52 -649 124
rect -615 -52 -609 124
rect -655 -64 -609 -52
rect -497 124 -451 136
rect -497 -52 -491 124
rect -457 -52 -451 124
rect -497 -64 -451 -52
rect -339 124 -293 136
rect -339 -52 -333 124
rect -299 -52 -293 124
rect -339 -64 -293 -52
rect -181 124 -135 136
rect -181 -52 -175 124
rect -141 -52 -135 124
rect -181 -64 -135 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 135 124 181 136
rect 135 -52 141 124
rect 175 -52 181 124
rect 135 -64 181 -52
rect 293 124 339 136
rect 293 -52 299 124
rect 333 -52 339 124
rect 293 -64 339 -52
rect 451 124 497 136
rect 451 -52 457 124
rect 491 -52 497 124
rect 451 -64 497 -52
rect 609 124 655 136
rect 609 -52 615 124
rect 649 -52 655 124
rect 609 -64 655 -52
rect 767 124 813 136
rect 767 -52 773 124
rect 807 -52 813 124
rect 767 -64 813 -52
rect 925 124 971 136
rect 925 -52 931 124
rect 965 -52 971 124
rect 925 -64 971 -52
rect 1083 124 1129 136
rect 1083 -52 1089 124
rect 1123 -52 1129 124
rect 1083 -64 1129 -52
rect 1241 124 1287 136
rect 1241 -52 1247 124
rect 1281 -52 1287 124
rect 1241 -64 1287 -52
rect 1399 124 1445 136
rect 1399 -52 1405 124
rect 1439 -52 1445 124
rect 1399 -64 1445 -52
rect 1557 124 1603 136
rect 1557 -52 1563 124
rect 1597 -52 1603 124
rect 1557 -64 1603 -52
rect -1547 -111 -1455 -105
rect -1547 -145 -1535 -111
rect -1467 -145 -1455 -111
rect -1547 -151 -1455 -145
rect -1389 -111 -1297 -105
rect -1389 -145 -1377 -111
rect -1309 -145 -1297 -111
rect -1389 -151 -1297 -145
rect -1231 -111 -1139 -105
rect -1231 -145 -1219 -111
rect -1151 -145 -1139 -111
rect -1231 -151 -1139 -145
rect -1073 -111 -981 -105
rect -1073 -145 -1061 -111
rect -993 -145 -981 -111
rect -1073 -151 -981 -145
rect -915 -111 -823 -105
rect -915 -145 -903 -111
rect -835 -145 -823 -111
rect -915 -151 -823 -145
rect -757 -111 -665 -105
rect -757 -145 -745 -111
rect -677 -145 -665 -111
rect -757 -151 -665 -145
rect -599 -111 -507 -105
rect -599 -145 -587 -111
rect -519 -145 -507 -111
rect -599 -151 -507 -145
rect -441 -111 -349 -105
rect -441 -145 -429 -111
rect -361 -145 -349 -111
rect -441 -151 -349 -145
rect -283 -111 -191 -105
rect -283 -145 -271 -111
rect -203 -145 -191 -111
rect -283 -151 -191 -145
rect -125 -111 -33 -105
rect -125 -145 -113 -111
rect -45 -145 -33 -111
rect -125 -151 -33 -145
rect 33 -111 125 -105
rect 33 -145 45 -111
rect 113 -145 125 -111
rect 33 -151 125 -145
rect 191 -111 283 -105
rect 191 -145 203 -111
rect 271 -145 283 -111
rect 191 -151 283 -145
rect 349 -111 441 -105
rect 349 -145 361 -111
rect 429 -145 441 -111
rect 349 -151 441 -145
rect 507 -111 599 -105
rect 507 -145 519 -111
rect 587 -145 599 -111
rect 507 -151 599 -145
rect 665 -111 757 -105
rect 665 -145 677 -111
rect 745 -145 757 -111
rect 665 -151 757 -145
rect 823 -111 915 -105
rect 823 -145 835 -111
rect 903 -145 915 -111
rect 823 -151 915 -145
rect 981 -111 1073 -105
rect 981 -145 993 -111
rect 1061 -145 1073 -111
rect 981 -151 1073 -145
rect 1139 -111 1231 -105
rect 1139 -145 1151 -111
rect 1219 -145 1231 -111
rect 1139 -151 1231 -145
rect 1297 -111 1389 -105
rect 1297 -145 1309 -111
rect 1377 -145 1389 -111
rect 1297 -151 1389 -145
rect 1455 -111 1547 -105
rect 1455 -145 1467 -111
rect 1535 -145 1547 -111
rect 1455 -151 1547 -145
<< labels >>
rlabel mvnsubdiffcont 0 -267 0 -267 0 B
port 1 nsew
rlabel mvpdiffc -1580 36 -1580 36 0 D0
port 2 nsew
rlabel polycont -1501 -128 -1501 -128 0 G0
port 3 nsew
rlabel mvpdiffc -1422 36 -1422 36 0 S1
port 4 nsew
rlabel polycont -1343 -128 -1343 -128 0 G1
port 5 nsew
rlabel mvpdiffc -1264 36 -1264 36 0 D2
port 6 nsew
rlabel polycont -1185 -128 -1185 -128 0 G2
port 7 nsew
rlabel mvpdiffc -1106 36 -1106 36 0 S3
port 8 nsew
rlabel polycont -1027 -128 -1027 -128 0 G3
port 9 nsew
rlabel mvpdiffc -948 36 -948 36 0 D4
port 10 nsew
rlabel polycont -869 -128 -869 -128 0 G4
port 11 nsew
rlabel mvpdiffc -790 36 -790 36 0 S5
port 12 nsew
rlabel polycont -711 -128 -711 -128 0 G5
port 13 nsew
rlabel mvpdiffc -632 36 -632 36 0 D6
port 14 nsew
rlabel polycont -553 -128 -553 -128 0 G6
port 15 nsew
rlabel mvpdiffc -474 36 -474 36 0 S7
port 16 nsew
rlabel polycont -395 -128 -395 -128 0 G7
port 17 nsew
rlabel mvpdiffc -316 36 -316 36 0 D8
port 18 nsew
rlabel polycont -237 -128 -237 -128 0 G8
port 19 nsew
rlabel mvpdiffc -158 36 -158 36 0 S9
port 20 nsew
rlabel polycont -79 -128 -79 -128 0 G9
port 21 nsew
rlabel mvpdiffc 0 36 0 36 0 D10
port 22 nsew
rlabel polycont 79 -128 79 -128 0 G10
port 23 nsew
rlabel mvpdiffc 158 36 158 36 0 S11
port 24 nsew
rlabel polycont 237 -128 237 -128 0 G11
port 25 nsew
rlabel mvpdiffc 316 36 316 36 0 D12
port 26 nsew
rlabel polycont 395 -128 395 -128 0 G12
port 27 nsew
rlabel mvpdiffc 474 36 474 36 0 S13
port 28 nsew
rlabel polycont 553 -128 553 -128 0 G13
port 29 nsew
rlabel mvpdiffc 632 36 632 36 0 D14
port 30 nsew
rlabel polycont 711 -128 711 -128 0 G14
port 31 nsew
rlabel mvpdiffc 790 36 790 36 0 S15
port 32 nsew
rlabel polycont 869 -128 869 -128 0 G15
port 33 nsew
rlabel mvpdiffc 948 36 948 36 0 D16
port 34 nsew
rlabel polycont 1027 -128 1027 -128 0 G16
port 35 nsew
rlabel mvpdiffc 1106 36 1106 36 0 S17
port 36 nsew
rlabel polycont 1185 -128 1185 -128 0 G17
port 37 nsew
rlabel mvpdiffc 1264 36 1264 36 0 D18
port 38 nsew
rlabel polycont 1343 -128 1343 -128 0 G18
port 39 nsew
rlabel mvpdiffc 1422 36 1422 36 0 S19
port 40 nsew
rlabel polycont 1501 -128 1501 -128 0 G19
port 41 nsew
<< properties >>
string FIXED_BBOX -1714 -267 1714 267
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
