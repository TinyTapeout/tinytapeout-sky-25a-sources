magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -236 -769 236 769
<< nmos >>
rect -50 -569 50 631
<< ndiff >>
rect -108 592 -50 631
rect -108 558 -96 592
rect -62 558 -50 592
rect -108 524 -50 558
rect -108 490 -96 524
rect -62 490 -50 524
rect -108 456 -50 490
rect -108 422 -96 456
rect -62 422 -50 456
rect -108 388 -50 422
rect -108 354 -96 388
rect -62 354 -50 388
rect -108 320 -50 354
rect -108 286 -96 320
rect -62 286 -50 320
rect -108 252 -50 286
rect -108 218 -96 252
rect -62 218 -50 252
rect -108 184 -50 218
rect -108 150 -96 184
rect -62 150 -50 184
rect -108 116 -50 150
rect -108 82 -96 116
rect -62 82 -50 116
rect -108 48 -50 82
rect -108 14 -96 48
rect -62 14 -50 48
rect -108 -20 -50 14
rect -108 -54 -96 -20
rect -62 -54 -50 -20
rect -108 -88 -50 -54
rect -108 -122 -96 -88
rect -62 -122 -50 -88
rect -108 -156 -50 -122
rect -108 -190 -96 -156
rect -62 -190 -50 -156
rect -108 -224 -50 -190
rect -108 -258 -96 -224
rect -62 -258 -50 -224
rect -108 -292 -50 -258
rect -108 -326 -96 -292
rect -62 -326 -50 -292
rect -108 -360 -50 -326
rect -108 -394 -96 -360
rect -62 -394 -50 -360
rect -108 -428 -50 -394
rect -108 -462 -96 -428
rect -62 -462 -50 -428
rect -108 -496 -50 -462
rect -108 -530 -96 -496
rect -62 -530 -50 -496
rect -108 -569 -50 -530
rect 50 592 108 631
rect 50 558 62 592
rect 96 558 108 592
rect 50 524 108 558
rect 50 490 62 524
rect 96 490 108 524
rect 50 456 108 490
rect 50 422 62 456
rect 96 422 108 456
rect 50 388 108 422
rect 50 354 62 388
rect 96 354 108 388
rect 50 320 108 354
rect 50 286 62 320
rect 96 286 108 320
rect 50 252 108 286
rect 50 218 62 252
rect 96 218 108 252
rect 50 184 108 218
rect 50 150 62 184
rect 96 150 108 184
rect 50 116 108 150
rect 50 82 62 116
rect 96 82 108 116
rect 50 48 108 82
rect 50 14 62 48
rect 96 14 108 48
rect 50 -20 108 14
rect 50 -54 62 -20
rect 96 -54 108 -20
rect 50 -88 108 -54
rect 50 -122 62 -88
rect 96 -122 108 -88
rect 50 -156 108 -122
rect 50 -190 62 -156
rect 96 -190 108 -156
rect 50 -224 108 -190
rect 50 -258 62 -224
rect 96 -258 108 -224
rect 50 -292 108 -258
rect 50 -326 62 -292
rect 96 -326 108 -292
rect 50 -360 108 -326
rect 50 -394 62 -360
rect 96 -394 108 -360
rect 50 -428 108 -394
rect 50 -462 62 -428
rect 96 -462 108 -428
rect 50 -496 108 -462
rect 50 -530 62 -496
rect 96 -530 108 -496
rect 50 -569 108 -530
<< ndiffc >>
rect -96 558 -62 592
rect -96 490 -62 524
rect -96 422 -62 456
rect -96 354 -62 388
rect -96 286 -62 320
rect -96 218 -62 252
rect -96 150 -62 184
rect -96 82 -62 116
rect -96 14 -62 48
rect -96 -54 -62 -20
rect -96 -122 -62 -88
rect -96 -190 -62 -156
rect -96 -258 -62 -224
rect -96 -326 -62 -292
rect -96 -394 -62 -360
rect -96 -462 -62 -428
rect -96 -530 -62 -496
rect 62 558 96 592
rect 62 490 96 524
rect 62 422 96 456
rect 62 354 96 388
rect 62 286 96 320
rect 62 218 96 252
rect 62 150 96 184
rect 62 82 96 116
rect 62 14 96 48
rect 62 -54 96 -20
rect 62 -122 96 -88
rect 62 -190 96 -156
rect 62 -258 96 -224
rect 62 -326 96 -292
rect 62 -394 96 -360
rect 62 -462 96 -428
rect 62 -530 96 -496
<< psubdiff >>
rect -210 709 -85 743
rect -51 709 -17 743
rect 17 709 51 743
rect 85 709 210 743
rect -210 629 -176 709
rect -210 561 -176 595
rect -210 493 -176 527
rect -210 425 -176 459
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -210 -459 -176 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect 176 629 210 709
rect 176 561 210 595
rect 176 493 210 527
rect 176 425 210 459
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect 176 -459 210 -425
rect 176 -527 210 -493
rect -210 -709 -176 -629
rect 176 -595 210 -561
rect 176 -709 210 -629
rect -210 -743 -85 -709
rect -51 -743 -17 -709
rect 17 -743 51 -709
rect 85 -743 210 -709
<< psubdiffcont >>
rect -85 709 -51 743
rect -17 709 17 743
rect 51 709 85 743
rect -210 595 -176 629
rect -210 527 -176 561
rect -210 459 -176 493
rect -210 391 -176 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect -210 -425 -176 -391
rect -210 -493 -176 -459
rect -210 -561 -176 -527
rect 176 595 210 629
rect 176 527 210 561
rect 176 459 210 493
rect 176 391 210 425
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect 176 -425 210 -391
rect 176 -493 210 -459
rect 176 -561 210 -527
rect -210 -629 -176 -595
rect 176 -629 210 -595
rect -85 -743 -51 -709
rect -17 -743 17 -709
rect 51 -743 85 -709
<< poly >>
rect -50 631 50 657
rect -50 -607 50 -569
rect -50 -641 -17 -607
rect 17 -641 50 -607
rect -50 -657 50 -641
<< polycont >>
rect -17 -641 17 -607
<< locali >>
rect -210 709 -85 743
rect -51 709 -17 743
rect 17 709 51 743
rect 85 709 210 743
rect -210 629 -176 709
rect -210 561 -176 595
rect -210 493 -176 527
rect -210 425 -176 459
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -210 -459 -176 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -96 592 -62 635
rect -96 524 -62 554
rect -96 456 -62 482
rect -96 388 -62 410
rect -96 320 -62 338
rect -96 252 -62 266
rect -96 184 -62 194
rect -96 116 -62 122
rect -96 48 -62 50
rect -96 12 -62 14
rect -96 -60 -62 -54
rect -96 -132 -62 -122
rect -96 -204 -62 -190
rect -96 -276 -62 -258
rect -96 -348 -62 -326
rect -96 -420 -62 -394
rect -96 -492 -62 -462
rect -96 -573 -62 -530
rect 62 592 96 635
rect 62 524 96 554
rect 62 456 96 482
rect 62 388 96 410
rect 62 320 96 338
rect 62 252 96 266
rect 62 184 96 194
rect 62 116 96 122
rect 62 48 96 50
rect 62 12 96 14
rect 62 -60 96 -54
rect 62 -132 96 -122
rect 62 -204 96 -190
rect 62 -276 96 -258
rect 62 -348 96 -326
rect 62 -420 96 -394
rect 62 -492 96 -462
rect 62 -573 96 -530
rect 176 629 210 709
rect 176 561 210 595
rect 176 493 210 527
rect 176 425 210 459
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect 176 -459 210 -425
rect 176 -527 210 -493
rect 176 -595 210 -561
rect -210 -709 -176 -629
rect -50 -641 -17 -607
rect 17 -641 50 -607
rect 176 -709 210 -629
rect -210 -743 -85 -709
rect -51 -743 -17 -709
rect 17 -743 51 -709
rect 85 -743 210 -709
<< viali >>
rect -96 558 -62 588
rect -96 554 -62 558
rect -96 490 -62 516
rect -96 482 -62 490
rect -96 422 -62 444
rect -96 410 -62 422
rect -96 354 -62 372
rect -96 338 -62 354
rect -96 286 -62 300
rect -96 266 -62 286
rect -96 218 -62 228
rect -96 194 -62 218
rect -96 150 -62 156
rect -96 122 -62 150
rect -96 82 -62 84
rect -96 50 -62 82
rect -96 -20 -62 12
rect -96 -22 -62 -20
rect -96 -88 -62 -60
rect -96 -94 -62 -88
rect -96 -156 -62 -132
rect -96 -166 -62 -156
rect -96 -224 -62 -204
rect -96 -238 -62 -224
rect -96 -292 -62 -276
rect -96 -310 -62 -292
rect -96 -360 -62 -348
rect -96 -382 -62 -360
rect -96 -428 -62 -420
rect -96 -454 -62 -428
rect -96 -496 -62 -492
rect -96 -526 -62 -496
rect 62 558 96 588
rect 62 554 96 558
rect 62 490 96 516
rect 62 482 96 490
rect 62 422 96 444
rect 62 410 96 422
rect 62 354 96 372
rect 62 338 96 354
rect 62 286 96 300
rect 62 266 96 286
rect 62 218 96 228
rect 62 194 96 218
rect 62 150 96 156
rect 62 122 96 150
rect 62 82 96 84
rect 62 50 96 82
rect 62 -20 96 12
rect 62 -22 96 -20
rect 62 -88 96 -60
rect 62 -94 96 -88
rect 62 -156 96 -132
rect 62 -166 96 -156
rect 62 -224 96 -204
rect 62 -238 96 -224
rect 62 -292 96 -276
rect 62 -310 96 -292
rect 62 -360 96 -348
rect 62 -382 96 -360
rect 62 -428 96 -420
rect 62 -454 96 -428
rect 62 -496 96 -492
rect 62 -526 96 -496
rect -17 -641 17 -607
<< metal1 >>
rect -102 588 -56 631
rect -102 554 -96 588
rect -62 554 -56 588
rect -102 516 -56 554
rect -102 482 -96 516
rect -62 482 -56 516
rect -102 444 -56 482
rect -102 410 -96 444
rect -62 410 -56 444
rect -102 372 -56 410
rect -102 338 -96 372
rect -62 338 -56 372
rect -102 300 -56 338
rect -102 266 -96 300
rect -62 266 -56 300
rect -102 228 -56 266
rect -102 194 -96 228
rect -62 194 -56 228
rect -102 156 -56 194
rect -102 122 -96 156
rect -62 122 -56 156
rect -102 84 -56 122
rect -102 50 -96 84
rect -62 50 -56 84
rect -102 12 -56 50
rect -102 -22 -96 12
rect -62 -22 -56 12
rect -102 -60 -56 -22
rect -102 -94 -96 -60
rect -62 -94 -56 -60
rect -102 -132 -56 -94
rect -102 -166 -96 -132
rect -62 -166 -56 -132
rect -102 -204 -56 -166
rect -102 -238 -96 -204
rect -62 -238 -56 -204
rect -102 -276 -56 -238
rect -102 -310 -96 -276
rect -62 -310 -56 -276
rect -102 -348 -56 -310
rect -102 -382 -96 -348
rect -62 -382 -56 -348
rect -102 -420 -56 -382
rect -102 -454 -96 -420
rect -62 -454 -56 -420
rect -102 -492 -56 -454
rect -102 -526 -96 -492
rect -62 -526 -56 -492
rect -102 -569 -56 -526
rect 56 588 102 631
rect 56 554 62 588
rect 96 554 102 588
rect 56 516 102 554
rect 56 482 62 516
rect 96 482 102 516
rect 56 444 102 482
rect 56 410 62 444
rect 96 410 102 444
rect 56 372 102 410
rect 56 338 62 372
rect 96 338 102 372
rect 56 300 102 338
rect 56 266 62 300
rect 96 266 102 300
rect 56 228 102 266
rect 56 194 62 228
rect 96 194 102 228
rect 56 156 102 194
rect 56 122 62 156
rect 96 122 102 156
rect 56 84 102 122
rect 56 50 62 84
rect 96 50 102 84
rect 56 12 102 50
rect 56 -22 62 12
rect 96 -22 102 12
rect 56 -60 102 -22
rect 56 -94 62 -60
rect 96 -94 102 -60
rect 56 -132 102 -94
rect 56 -166 62 -132
rect 96 -166 102 -132
rect 56 -204 102 -166
rect 56 -238 62 -204
rect 96 -238 102 -204
rect 56 -276 102 -238
rect 56 -310 62 -276
rect 96 -310 102 -276
rect 56 -348 102 -310
rect 56 -382 62 -348
rect 96 -382 102 -348
rect 56 -420 102 -382
rect 56 -454 62 -420
rect 96 -454 102 -420
rect 56 -492 102 -454
rect 56 -526 62 -492
rect 96 -526 102 -492
rect 56 -569 102 -526
rect -46 -607 46 -601
rect -46 -641 -17 -607
rect 17 -641 46 -607
rect -46 -647 46 -641
<< properties >>
string FIXED_BBOX -193 -726 193 726
<< end >>
