magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 704 240
<< ptap >>
rect -48 60 752 100
rect -48 100 752 140
rect -48 140 752 180
rect -48 180 48 220
rect 656 180 752 220
rect -48 220 48 260
rect 656 220 752 260
<< locali >>
rect -48 60 752 100
rect -48 100 752 140
rect -48 140 752 180
rect -48 180 48 220
rect 656 180 752 220
rect -48 220 48 260
rect 656 220 752 260
<< ptapc >>
rect 80 100 592 140
<< pwell >>
rect -92 -64 796 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 704 240
<< end >>
