magic
tech sky130A
magscale 1 2
timestamp 1752660100
<< nwell >>
rect -936 -2332 946 2342
<< pmoslvt >>
rect -740 123 -540 2123
rect -482 123 -282 2123
rect -224 123 -24 2123
rect 34 123 234 2123
rect 292 123 492 2123
rect 550 123 750 2123
rect -740 -2113 -540 -113
rect -482 -2113 -282 -113
rect -224 -2113 -24 -113
rect 34 -2113 234 -113
rect 292 -2113 492 -113
rect 550 -2113 750 -113
<< pdiff >>
rect -798 2111 -740 2123
rect -798 135 -786 2111
rect -752 135 -740 2111
rect -798 123 -740 135
rect -540 2111 -482 2123
rect -540 135 -528 2111
rect -494 135 -482 2111
rect -540 123 -482 135
rect -282 2111 -224 2123
rect -282 135 -270 2111
rect -236 135 -224 2111
rect -282 123 -224 135
rect -24 2111 34 2123
rect -24 135 -12 2111
rect 22 135 34 2111
rect -24 123 34 135
rect 234 2111 292 2123
rect 234 135 246 2111
rect 280 135 292 2111
rect 234 123 292 135
rect 492 2111 550 2123
rect 492 135 504 2111
rect 538 135 550 2111
rect 492 123 550 135
rect 750 2111 808 2123
rect 750 135 762 2111
rect 796 135 808 2111
rect 750 123 808 135
rect -798 -125 -740 -113
rect -798 -2101 -786 -125
rect -752 -2101 -740 -125
rect -798 -2113 -740 -2101
rect -540 -125 -482 -113
rect -540 -2101 -528 -125
rect -494 -2101 -482 -125
rect -540 -2113 -482 -2101
rect -282 -125 -224 -113
rect -282 -2101 -270 -125
rect -236 -2101 -224 -125
rect -282 -2113 -224 -2101
rect -24 -125 34 -113
rect -24 -2101 -12 -125
rect 22 -2101 34 -125
rect -24 -2113 34 -2101
rect 234 -125 292 -113
rect 234 -2101 246 -125
rect 280 -2101 292 -125
rect 234 -2113 292 -2101
rect 492 -125 550 -113
rect 492 -2101 504 -125
rect 538 -2101 550 -125
rect 492 -2113 550 -2101
rect 750 -125 808 -113
rect 750 -2101 762 -125
rect 796 -2101 808 -125
rect 750 -2113 808 -2101
<< pdiffc >>
rect -786 135 -752 2111
rect -528 135 -494 2111
rect -270 135 -236 2111
rect -12 135 22 2111
rect 246 135 280 2111
rect 504 135 538 2111
rect 762 135 796 2111
rect -786 -2101 -752 -125
rect -528 -2101 -494 -125
rect -270 -2101 -236 -125
rect -12 -2101 22 -125
rect 246 -2101 280 -125
rect 504 -2101 538 -125
rect 762 -2101 796 -125
<< nsubdiff >>
rect -900 2272 -804 2306
rect 814 2272 910 2306
rect -900 2210 -866 2272
rect 876 2210 910 2272
rect -900 -2262 -866 -2200
rect 876 -2262 910 -2200
rect -900 -2296 -804 -2262
rect 814 -2296 910 -2262
<< nsubdiffcont >>
rect -804 2272 814 2306
rect -900 -2200 -866 2210
rect 876 -2200 910 2210
rect -804 -2296 814 -2262
<< poly >>
rect -740 2204 -540 2220
rect -740 2170 -724 2204
rect -556 2170 -540 2204
rect -740 2123 -540 2170
rect -482 2204 -282 2220
rect -482 2170 -466 2204
rect -298 2170 -282 2204
rect -482 2123 -282 2170
rect -224 2204 -24 2220
rect -224 2170 -208 2204
rect -40 2170 -24 2204
rect -224 2123 -24 2170
rect 34 2204 234 2220
rect 34 2170 50 2204
rect 218 2170 234 2204
rect 34 2123 234 2170
rect 292 2204 492 2220
rect 292 2170 308 2204
rect 476 2170 492 2204
rect 292 2123 492 2170
rect 550 2204 750 2220
rect 550 2170 566 2204
rect 734 2170 750 2204
rect 550 2123 750 2170
rect -740 76 -540 123
rect -740 42 -724 76
rect -556 42 -540 76
rect -740 26 -540 42
rect -482 76 -282 123
rect -482 42 -466 76
rect -298 42 -282 76
rect -482 26 -282 42
rect -224 76 -24 123
rect -224 42 -208 76
rect -40 42 -24 76
rect -224 26 -24 42
rect 34 76 234 123
rect 34 42 50 76
rect 218 42 234 76
rect 34 26 234 42
rect 292 76 492 123
rect 292 42 308 76
rect 476 42 492 76
rect 292 26 492 42
rect 550 76 750 123
rect 550 42 566 76
rect 734 42 750 76
rect 550 26 750 42
rect -740 -32 -540 -16
rect -740 -66 -724 -32
rect -556 -66 -540 -32
rect -740 -113 -540 -66
rect -482 -32 -282 -16
rect -482 -66 -466 -32
rect -298 -66 -282 -32
rect -482 -113 -282 -66
rect -224 -32 -24 -16
rect -224 -66 -208 -32
rect -40 -66 -24 -32
rect -224 -113 -24 -66
rect 34 -32 234 -16
rect 34 -66 50 -32
rect 218 -66 234 -32
rect 34 -113 234 -66
rect 292 -32 492 -16
rect 292 -66 308 -32
rect 476 -66 492 -32
rect 292 -113 492 -66
rect 550 -32 750 -16
rect 550 -66 566 -32
rect 734 -66 750 -32
rect 550 -113 750 -66
rect -740 -2160 -540 -2113
rect -740 -2194 -724 -2160
rect -556 -2194 -540 -2160
rect -740 -2210 -540 -2194
rect -482 -2160 -282 -2113
rect -482 -2194 -466 -2160
rect -298 -2194 -282 -2160
rect -482 -2210 -282 -2194
rect -224 -2160 -24 -2113
rect -224 -2194 -208 -2160
rect -40 -2194 -24 -2160
rect -224 -2210 -24 -2194
rect 34 -2160 234 -2113
rect 34 -2194 50 -2160
rect 218 -2194 234 -2160
rect 34 -2210 234 -2194
rect 292 -2160 492 -2113
rect 292 -2194 308 -2160
rect 476 -2194 492 -2160
rect 292 -2210 492 -2194
rect 550 -2160 750 -2113
rect 550 -2194 566 -2160
rect 734 -2194 750 -2160
rect 550 -2210 750 -2194
<< polycont >>
rect -724 2170 -556 2204
rect -466 2170 -298 2204
rect -208 2170 -40 2204
rect 50 2170 218 2204
rect 308 2170 476 2204
rect 566 2170 734 2204
rect -724 42 -556 76
rect -466 42 -298 76
rect -208 42 -40 76
rect 50 42 218 76
rect 308 42 476 76
rect 566 42 734 76
rect -724 -66 -556 -32
rect -466 -66 -298 -32
rect -208 -66 -40 -32
rect 50 -66 218 -32
rect 308 -66 476 -32
rect 566 -66 734 -32
rect -724 -2194 -556 -2160
rect -466 -2194 -298 -2160
rect -208 -2194 -40 -2160
rect 50 -2194 218 -2160
rect 308 -2194 476 -2160
rect 566 -2194 734 -2160
<< locali >>
rect -900 2272 -804 2306
rect 814 2272 910 2306
rect -900 2210 -866 2272
rect 876 2210 910 2272
rect -740 2170 -724 2204
rect -556 2170 -540 2204
rect -482 2170 -466 2204
rect -298 2170 -282 2204
rect -224 2170 -208 2204
rect -40 2170 -24 2204
rect 34 2170 50 2204
rect 218 2170 234 2204
rect 292 2170 308 2204
rect 476 2170 492 2204
rect 550 2170 566 2204
rect 734 2170 750 2204
rect -786 2111 -752 2127
rect -786 119 -752 135
rect -528 2111 -494 2127
rect -528 119 -494 135
rect -270 2111 -236 2127
rect -270 119 -236 135
rect -12 2111 22 2127
rect -12 119 22 135
rect 246 2111 280 2127
rect 246 119 280 135
rect 504 2111 538 2127
rect 504 119 538 135
rect 762 2111 796 2127
rect 762 119 796 135
rect -740 42 -724 76
rect -556 42 -540 76
rect -482 42 -466 76
rect -298 42 -282 76
rect -224 42 -208 76
rect -40 42 -24 76
rect 34 42 50 76
rect 218 42 234 76
rect 292 42 308 76
rect 476 42 492 76
rect 550 42 566 76
rect 734 42 750 76
rect -740 -66 -724 -32
rect -556 -66 -540 -32
rect -482 -66 -466 -32
rect -298 -66 -282 -32
rect -224 -66 -208 -32
rect -40 -66 -24 -32
rect 34 -66 50 -32
rect 218 -66 234 -32
rect 292 -66 308 -32
rect 476 -66 492 -32
rect 550 -66 566 -32
rect 734 -66 750 -32
rect -786 -125 -752 -109
rect -786 -2117 -752 -2101
rect -528 -125 -494 -109
rect -528 -2117 -494 -2101
rect -270 -125 -236 -109
rect -270 -2117 -236 -2101
rect -12 -125 22 -109
rect -12 -2117 22 -2101
rect 246 -125 280 -109
rect 246 -2117 280 -2101
rect 504 -125 538 -109
rect 504 -2117 538 -2101
rect 762 -125 796 -109
rect 762 -2117 796 -2101
rect -740 -2194 -724 -2160
rect -556 -2194 -540 -2160
rect -482 -2194 -466 -2160
rect -298 -2194 -282 -2160
rect -224 -2194 -208 -2160
rect -40 -2194 -24 -2160
rect 34 -2194 50 -2160
rect 218 -2194 234 -2160
rect 292 -2194 308 -2160
rect 476 -2194 492 -2160
rect 550 -2194 566 -2160
rect 734 -2194 750 -2160
rect -900 -2262 -866 -2200
rect 876 -2262 910 -2200
rect -900 -2296 -804 -2262
rect 814 -2296 910 -2262
<< viali >>
rect -724 2170 -556 2204
rect -466 2170 -298 2204
rect -208 2170 -40 2204
rect 50 2170 218 2204
rect 308 2170 476 2204
rect 566 2170 734 2204
rect -786 135 -752 2111
rect -528 135 -494 2111
rect -270 135 -236 2111
rect -12 135 22 2111
rect 246 135 280 2111
rect 504 135 538 2111
rect 762 135 796 2111
rect -724 42 -556 76
rect -466 42 -298 76
rect -208 42 -40 76
rect 50 42 218 76
rect 308 42 476 76
rect 566 42 734 76
rect -724 -66 -556 -32
rect -466 -66 -298 -32
rect -208 -66 -40 -32
rect 50 -66 218 -32
rect 308 -66 476 -32
rect 566 -66 734 -32
rect -786 -2101 -752 -125
rect -528 -2101 -494 -125
rect -270 -2101 -236 -125
rect -12 -2101 22 -125
rect 246 -2101 280 -125
rect 504 -2101 538 -125
rect 762 -2101 796 -125
rect -724 -2194 -556 -2160
rect -466 -2194 -298 -2160
rect -208 -2194 -40 -2160
rect 50 -2194 218 -2160
rect 308 -2194 476 -2160
rect 566 -2194 734 -2160
<< metal1 >>
rect -736 2204 -544 2210
rect -736 2170 -724 2204
rect -556 2170 -544 2204
rect -736 2164 -544 2170
rect -478 2204 -286 2210
rect -478 2170 -466 2204
rect -298 2170 -286 2204
rect -478 2164 -286 2170
rect -220 2204 -28 2210
rect -220 2170 -208 2204
rect -40 2170 -28 2204
rect -220 2164 -28 2170
rect 38 2204 230 2210
rect 38 2170 50 2204
rect 218 2170 230 2204
rect 38 2164 230 2170
rect 296 2204 488 2210
rect 296 2170 308 2204
rect 476 2170 488 2204
rect 296 2164 488 2170
rect 554 2204 746 2210
rect 554 2170 566 2204
rect 734 2170 746 2204
rect 554 2164 746 2170
rect -792 2111 -746 2123
rect -792 135 -786 2111
rect -752 135 -746 2111
rect -792 123 -746 135
rect -534 2111 -488 2123
rect -534 135 -528 2111
rect -494 135 -488 2111
rect -534 123 -488 135
rect -276 2111 -230 2123
rect -276 135 -270 2111
rect -236 135 -230 2111
rect -276 123 -230 135
rect -18 2111 28 2123
rect -18 135 -12 2111
rect 22 135 28 2111
rect -18 123 28 135
rect 240 2111 286 2123
rect 240 135 246 2111
rect 280 135 286 2111
rect 240 123 286 135
rect 498 2111 544 2123
rect 498 135 504 2111
rect 538 135 544 2111
rect 498 123 544 135
rect 756 2111 802 2123
rect 756 135 762 2111
rect 796 135 802 2111
rect 756 123 802 135
rect -736 76 -544 82
rect -736 42 -724 76
rect -556 42 -544 76
rect -736 36 -544 42
rect -478 76 -286 82
rect -478 42 -466 76
rect -298 42 -286 76
rect -478 36 -286 42
rect -220 76 -28 82
rect -220 42 -208 76
rect -40 42 -28 76
rect -220 36 -28 42
rect 38 76 230 82
rect 38 42 50 76
rect 218 42 230 76
rect 38 36 230 42
rect 296 76 488 82
rect 296 42 308 76
rect 476 42 488 76
rect 296 36 488 42
rect 554 76 746 82
rect 554 42 566 76
rect 734 42 746 76
rect 554 36 746 42
rect -736 -32 -544 -26
rect -736 -66 -724 -32
rect -556 -66 -544 -32
rect -736 -72 -544 -66
rect -478 -32 -286 -26
rect -478 -66 -466 -32
rect -298 -66 -286 -32
rect -478 -72 -286 -66
rect -220 -32 -28 -26
rect -220 -66 -208 -32
rect -40 -66 -28 -32
rect -220 -72 -28 -66
rect 38 -32 230 -26
rect 38 -66 50 -32
rect 218 -66 230 -32
rect 38 -72 230 -66
rect 296 -32 488 -26
rect 296 -66 308 -32
rect 476 -66 488 -32
rect 296 -72 488 -66
rect 554 -32 746 -26
rect 554 -66 566 -32
rect 734 -66 746 -32
rect 554 -72 746 -66
rect -792 -125 -746 -113
rect -792 -2101 -786 -125
rect -752 -2101 -746 -125
rect -792 -2113 -746 -2101
rect -534 -125 -488 -113
rect -534 -2101 -528 -125
rect -494 -2101 -488 -125
rect -534 -2113 -488 -2101
rect -276 -125 -230 -113
rect -276 -2101 -270 -125
rect -236 -2101 -230 -125
rect -276 -2113 -230 -2101
rect -18 -125 28 -113
rect -18 -2101 -12 -125
rect 22 -2101 28 -125
rect -18 -2113 28 -2101
rect 240 -125 286 -113
rect 240 -2101 246 -125
rect 280 -2101 286 -125
rect 240 -2113 286 -2101
rect 498 -125 544 -113
rect 498 -2101 504 -125
rect 538 -2101 544 -125
rect 498 -2113 544 -2101
rect 756 -125 802 -113
rect 756 -2101 762 -125
rect 796 -2101 802 -125
rect 756 -2113 802 -2101
rect -736 -2160 -544 -2154
rect -736 -2194 -724 -2160
rect -556 -2194 -544 -2160
rect -736 -2200 -544 -2194
rect -478 -2160 -286 -2154
rect -478 -2194 -466 -2160
rect -298 -2194 -286 -2160
rect -478 -2200 -286 -2194
rect -220 -2160 -28 -2154
rect -220 -2194 -208 -2160
rect -40 -2194 -28 -2160
rect -220 -2200 -28 -2194
rect 38 -2160 230 -2154
rect 38 -2194 50 -2160
rect 218 -2194 230 -2160
rect 38 -2200 230 -2194
rect 296 -2160 488 -2154
rect 296 -2194 308 -2160
rect 476 -2194 488 -2160
rect 296 -2200 488 -2194
rect 554 -2160 746 -2154
rect 554 -2194 566 -2160
rect 734 -2194 746 -2160
rect 554 -2200 746 -2194
<< properties >>
string FIXED_BBOX -883 -2279 893 2289
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
