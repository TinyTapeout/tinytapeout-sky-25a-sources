// Generated from: 20250914-213301_binTestAcc9744_seed445809_epochs100_2x2560_b256_lr50_interconnect.npz

module net (
    input  wire [254:0] in,
    output wire [2559:0] out,
    output wire [2549:0] categories
);
    wire [2560:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = ~(in[9] ^ in[36]); 
    assign layer_0[1] = in[230] | in[119]; 
    assign layer_0[2] = in[106] | in[66]; 
    assign layer_0[3] = ~in[137] | (in[90] & in[137]); 
    assign layer_0[4] = in[59] ^ in[39]; 
    assign layer_0[5] = ~(in[249] ^ in[246]); 
    assign layer_0[6] = in[9] & ~in[76]; 
    assign layer_0[7] = ~in[54] | (in[24] & in[54]); 
    assign layer_0[8] = ~(in[141] ^ in[175]); 
    assign layer_0[9] = in[151] ^ in[120]; 
    assign layer_0[10] = in[124] ^ in[106]; 
    assign layer_0[11] = ~(in[194] | in[123]); 
    assign layer_0[12] = in[168] | in[51]; 
    assign layer_0[13] = ~(in[162] | in[163]); 
    assign layer_0[14] = in[95] & ~in[139]; 
    assign layer_0[15] = in[236] ^ in[249]; 
    assign layer_0[16] = ~in[75] | (in[232] & in[75]); 
    assign layer_0[17] = in[186] & ~in[95]; 
    assign layer_0[18] = ~(in[60] | in[75]); 
    assign layer_0[19] = in[201] | in[203]; 
    assign layer_0[20] = in[104] ^ in[61]; 
    assign layer_0[21] = ~(in[210] ^ in[231]); 
    assign layer_0[22] = in[196] ^ in[227]; 
    assign layer_0[23] = in[102] | in[47]; 
    assign layer_0[24] = in[116] ^ in[114]; 
    assign layer_0[25] = in[242] ^ in[185]; 
    assign layer_0[26] = ~(in[149] ^ in[163]); 
    assign layer_0[27] = in[40] | in[56]; 
    assign layer_0[28] = in[40] ^ in[87]; 
    assign layer_0[29] = ~in[188] | (in[91] & in[188]); 
    assign layer_0[30] = in[104] & ~in[156]; 
    assign layer_0[31] = in[189] ^ in[107]; 
    assign layer_0[32] = ~(in[248] | in[104]); 
    assign layer_0[33] = ~(in[102] ^ in[155]); 
    assign layer_0[34] = in[228] & ~in[209]; 
    assign layer_0[35] = ~in[69] | (in[69] & in[66]); 
    assign layer_0[36] = ~(in[155] | in[92]); 
    assign layer_0[37] = ~(in[230] | in[215]); 
    assign layer_0[38] = ~(in[235] | in[60]); 
    assign layer_0[39] = in[130] | in[148]; 
    assign layer_0[40] = in[83] & ~in[118]; 
    assign layer_0[41] = ~(in[79] ^ in[46]); 
    assign layer_0[42] = 1'b1; 
    assign layer_0[43] = in[154]; 
    assign layer_0[44] = in[150]; 
    assign layer_0[45] = in[77] ^ in[78]; 
    assign layer_0[46] = ~in[197] | (in[79] & in[197]); 
    assign layer_0[47] = ~(in[172] | in[180]); 
    assign layer_0[48] = ~(in[244] ^ in[182]); 
    assign layer_0[49] = ~in[117]; 
    assign layer_0[50] = ~(in[130] ^ in[116]); 
    assign layer_0[51] = ~(in[166] ^ in[164]); 
    assign layer_0[52] = in[70] ^ in[101]; 
    assign layer_0[53] = ~in[193]; 
    assign layer_0[54] = in[25] | in[28]; 
    assign layer_0[55] = ~(in[218] ^ in[195]); 
    assign layer_0[56] = in[164] ^ in[229]; 
    assign layer_0[57] = in[246] | in[243]; 
    assign layer_0[58] = in[214] & ~in[123]; 
    assign layer_0[59] = ~in[170]; 
    assign layer_0[60] = in[138] ^ in[184]; 
    assign layer_0[61] = in[55] | in[140]; 
    assign layer_0[62] = ~(in[167] ^ in[88]); 
    assign layer_0[63] = ~(in[187] ^ in[249]); 
    assign layer_0[64] = ~(in[105] ^ in[90]); 
    assign layer_0[65] = ~in[114] | (in[101] & in[114]); 
    assign layer_0[66] = in[138] ^ in[185]; 
    assign layer_0[67] = ~(in[173] ^ in[221]); 
    assign layer_0[68] = in[185]; 
    assign layer_0[69] = ~in[137] | (in[193] & in[137]); 
    assign layer_0[70] = in[59] ^ in[119]; 
    assign layer_0[71] = in[87] ^ in[85]; 
    assign layer_0[72] = in[93] ^ in[216]; 
    assign layer_0[73] = ~(in[164] ^ in[146]); 
    assign layer_0[74] = ~(in[71] ^ in[73]); 
    assign layer_0[75] = in[193] | in[8]; 
    assign layer_0[76] = ~(in[175] ^ in[209]); 
    assign layer_0[77] = ~(in[11] | in[152]); 
    assign layer_0[78] = ~(in[230] | in[110]); 
    assign layer_0[79] = in[146] & ~in[89]; 
    assign layer_0[80] = ~in[185] | (in[214] & in[185]); 
    assign layer_0[81] = ~(in[102] ^ in[100]); 
    assign layer_0[82] = in[164] ^ in[132]; 
    assign layer_0[83] = ~(in[113] | in[138]); 
    assign layer_0[84] = in[88] & ~in[197]; 
    assign layer_0[85] = in[187] ^ in[196]; 
    assign layer_0[86] = ~in[78]; 
    assign layer_0[87] = ~in[54]; 
    assign layer_0[88] = ~in[137] | (in[137] & in[22]); 
    assign layer_0[89] = in[46] ^ in[63]; 
    assign layer_0[90] = in[69] ^ in[38]; 
    assign layer_0[91] = in[251] | in[219]; 
    assign layer_0[92] = in[149] | in[51]; 
    assign layer_0[93] = in[42] ^ in[73]; 
    assign layer_0[94] = in[250] ^ in[247]; 
    assign layer_0[95] = ~(in[188] ^ in[219]); 
    assign layer_0[96] = ~in[154] | (in[136] & in[154]); 
    assign layer_0[97] = ~(in[250] ^ in[233]); 
    assign layer_0[98] = ~(in[51] ^ in[202]); 
    assign layer_0[99] = ~(in[172] ^ in[174]); 
    assign layer_0[100] = in[145] & ~in[53]; 
    assign layer_0[101] = ~(in[195] | in[197]); 
    assign layer_0[102] = in[38] | in[137]; 
    assign layer_0[103] = ~(in[159] | in[11]); 
    assign layer_0[104] = in[6] ^ in[242]; 
    assign layer_0[105] = in[72] & ~in[167]; 
    assign layer_0[106] = ~(in[198] ^ in[167]); 
    assign layer_0[107] = in[183] ^ in[81]; 
    assign layer_0[108] = in[74]; 
    assign layer_0[109] = ~(in[122] ^ in[197]); 
    assign layer_0[110] = ~in[169]; 
    assign layer_0[111] = in[102] ^ in[39]; 
    assign layer_0[112] = in[211] | in[220]; 
    assign layer_0[113] = ~in[166]; 
    assign layer_0[114] = ~in[138]; 
    assign layer_0[115] = in[5] | in[9]; 
    assign layer_0[116] = in[3]; 
    assign layer_0[117] = ~(in[182] ^ in[180]); 
    assign layer_0[118] = in[235] ^ in[35]; 
    assign layer_0[119] = ~(in[107] ^ in[156]); 
    assign layer_0[120] = in[122]; 
    assign layer_0[121] = ~(in[184] ^ in[152]); 
    assign layer_0[122] = ~in[183] | (in[183] & in[89]); 
    assign layer_0[123] = ~(in[102] ^ in[115]); 
    assign layer_0[124] = ~in[215] | (in[123] & in[215]); 
    assign layer_0[125] = ~(in[72] ^ in[41]); 
    assign layer_0[126] = in[182] | in[146]; 
    assign layer_0[127] = in[234] | in[120]; 
    assign layer_0[128] = ~(in[26] ^ in[170]); 
    assign layer_0[129] = in[84] ^ in[98]; 
    assign layer_0[130] = ~(in[250] ^ in[236]); 
    assign layer_0[131] = ~in[169] | (in[169] & in[132]); 
    assign layer_0[132] = ~(in[199] | in[100]); 
    assign layer_0[133] = ~(in[180] ^ in[244]); 
    assign layer_0[134] = ~(in[121] ^ in[89]); 
    assign layer_0[135] = ~(in[138] | in[44]); 
    assign layer_0[136] = in[39] ^ in[71]; 
    assign layer_0[137] = in[58] ^ in[89]; 
    assign layer_0[138] = ~(in[117] ^ in[135]); 
    assign layer_0[139] = in[84] & in[130]; 
    assign layer_0[140] = in[84] ^ in[86]; 
    assign layer_0[141] = ~(in[46] ^ in[92]); 
    assign layer_0[142] = in[71] ^ in[38]; 
    assign layer_0[143] = ~(in[248] ^ in[250]); 
    assign layer_0[144] = in[88] | in[120]; 
    assign layer_0[145] = ~(in[132] ^ in[118]); 
    assign layer_0[146] = in[9] | in[130]; 
    assign layer_0[147] = in[233]; 
    assign layer_0[148] = in[154] & ~in[80]; 
    assign layer_0[149] = ~in[47]; 
    assign layer_0[150] = in[125] | in[114]; 
    assign layer_0[151] = ~(in[130] | in[131]); 
    assign layer_0[152] = in[77] | in[41]; 
    assign layer_0[153] = in[52] ^ in[155]; 
    assign layer_0[154] = ~(in[199] | in[230]); 
    assign layer_0[155] = in[131] ^ in[117]; 
    assign layer_0[156] = in[200] & ~in[41]; 
    assign layer_0[157] = ~(in[22] ^ in[214]); 
    assign layer_0[158] = in[94] | in[212]; 
    assign layer_0[159] = in[213] ^ in[211]; 
    assign layer_0[160] = ~(in[99] ^ in[101]); 
    assign layer_0[161] = ~(in[102] ^ in[70]); 
    assign layer_0[162] = ~in[57] | (in[57] & in[183]); 
    assign layer_0[163] = ~(in[104] | in[79]); 
    assign layer_0[164] = in[213] & ~in[123]; 
    assign layer_0[165] = ~(in[60] ^ in[88]); 
    assign layer_0[166] = in[94] ^ in[107]; 
    assign layer_0[167] = ~(in[91] | in[105]); 
    assign layer_0[168] = in[91] & ~in[27]; 
    assign layer_0[169] = ~in[125]; 
    assign layer_0[170] = ~in[72] | (in[63] & in[72]); 
    assign layer_0[171] = ~(in[82] ^ in[154]); 
    assign layer_0[172] = ~in[121]; 
    assign layer_0[173] = ~(in[167] | in[148]); 
    assign layer_0[174] = ~(in[142] | in[104]); 
    assign layer_0[175] = in[39] ^ in[123]; 
    assign layer_0[176] = in[185] ^ in[218]; 
    assign layer_0[177] = in[28] ^ in[124]; 
    assign layer_0[178] = in[11]; 
    assign layer_0[179] = in[134] ^ in[213]; 
    assign layer_0[180] = in[121]; 
    assign layer_0[181] = ~(in[167] ^ in[124]); 
    assign layer_0[182] = ~in[232] | (in[232] & in[149]); 
    assign layer_0[183] = in[109] ^ in[78]; 
    assign layer_0[184] = ~in[153] | (in[153] & in[5]); 
    assign layer_0[185] = ~(in[101] | in[217]); 
    assign layer_0[186] = in[35] | in[196]; 
    assign layer_0[187] = in[183] | in[20]; 
    assign layer_0[188] = ~(in[6] | in[8]); 
    assign layer_0[189] = in[76] ^ in[213]; 
    assign layer_0[190] = ~(in[11] ^ in[12]); 
    assign layer_0[191] = in[9] | in[137]; 
    assign layer_0[192] = in[116] & ~in[180]; 
    assign layer_0[193] = in[108] ^ in[90]; 
    assign layer_0[194] = ~(in[149] ^ in[132]); 
    assign layer_0[195] = in[42] | in[67]; 
    assign layer_0[196] = in[104] ^ in[90]; 
    assign layer_0[197] = ~(in[199] ^ in[69]); 
    assign layer_0[198] = ~(in[108] ^ in[78]); 
    assign layer_0[199] = ~(in[156] | in[139]); 
    assign layer_0[200] = in[130] ^ in[132]; 
    assign layer_0[201] = ~(in[117] ^ in[131]); 
    assign layer_0[202] = in[187] ^ in[218]; 
    assign layer_0[203] = ~(in[163] ^ in[100]); 
    assign layer_0[204] = in[229]; 
    assign layer_0[205] = ~(in[136] ^ in[167]); 
    assign layer_0[206] = in[5] | in[173]; 
    assign layer_0[207] = ~(in[124] | in[74]); 
    assign layer_0[208] = in[113] ^ in[115]; 
    assign layer_0[209] = in[120] ^ in[88]; 
    assign layer_0[210] = in[97] ^ in[84]; 
    assign layer_0[211] = ~(in[156] ^ in[138]); 
    assign layer_0[212] = ~(in[243] | in[105]); 
    assign layer_0[213] = ~in[137] | (in[137] & in[92]); 
    assign layer_0[214] = ~in[203]; 
    assign layer_0[215] = ~(in[139] ^ in[82]); 
    assign layer_0[216] = in[83] | in[69]; 
    assign layer_0[217] = in[184] | in[215]; 
    assign layer_0[218] = in[26] | in[135]; 
    assign layer_0[219] = in[156] | in[36]; 
    assign layer_0[220] = ~in[99]; 
    assign layer_0[221] = ~(in[37] ^ in[78]); 
    assign layer_0[222] = in[88] ^ in[119]; 
    assign layer_0[223] = in[141] | in[162]; 
    assign layer_0[224] = in[182]; 
    assign layer_0[225] = in[99]; 
    assign layer_0[226] = in[90] ^ in[194]; 
    assign layer_0[227] = in[171] ^ in[140]; 
    assign layer_0[228] = in[157] ^ in[86]; 
    assign layer_0[229] = in[104] ^ in[89]; 
    assign layer_0[230] = ~in[151]; 
    assign layer_0[231] = ~in[186]; 
    assign layer_0[232] = in[154] & in[185]; 
    assign layer_0[233] = in[117] | in[147]; 
    assign layer_0[234] = in[90] ^ in[108]; 
    assign layer_0[235] = ~(in[49] ^ in[158]); 
    assign layer_0[236] = ~(in[235] | in[199]); 
    assign layer_0[237] = ~(in[198] & in[151]); 
    assign layer_0[238] = ~(in[27] ^ in[24]); 
    assign layer_0[239] = ~(in[235] | in[204]); 
    assign layer_0[240] = in[122] & ~in[94]; 
    assign layer_0[241] = in[210] ^ in[245]; 
    assign layer_0[242] = ~(in[181] ^ in[85]); 
    assign layer_0[243] = ~in[141]; 
    assign layer_0[244] = in[87] ^ in[101]; 
    assign layer_0[245] = ~in[109]; 
    assign layer_0[246] = in[67] | in[69]; 
    assign layer_0[247] = ~(in[199] | in[214]); 
    assign layer_0[248] = in[158] | in[58]; 
    assign layer_0[249] = ~in[137] | (in[137] & in[184]); 
    assign layer_0[250] = ~(in[27] ^ in[142]); 
    assign layer_0[251] = ~(in[165] | in[182]); 
    assign layer_0[252] = ~(in[118] | in[172]); 
    assign layer_0[253] = ~(in[43] ^ in[74]); 
    assign layer_0[254] = in[51] & ~in[251]; 
    assign layer_0[255] = in[105] & ~in[9]; 
    assign layer_0[256] = in[60] | in[78]; 
    assign layer_0[257] = in[105] ^ in[113]; 
    assign layer_0[258] = ~(in[29] | in[190]); 
    assign layer_0[259] = in[126] | in[28]; 
    assign layer_0[260] = in[247] | in[231]; 
    assign layer_0[261] = in[155] | in[158]; 
    assign layer_0[262] = in[98] | in[110]; 
    assign layer_0[263] = ~in[6]; 
    assign layer_0[264] = in[43] ^ in[106]; 
    assign layer_0[265] = in[227] ^ in[72]; 
    assign layer_0[266] = in[209] ^ in[217]; 
    assign layer_0[267] = in[213]; 
    assign layer_0[268] = in[109] & ~in[249]; 
    assign layer_0[269] = ~in[86] | (in[86] & in[21]); 
    assign layer_0[270] = ~(in[89] | in[231]); 
    assign layer_0[271] = ~(in[229] | in[189]); 
    assign layer_0[272] = in[168] | in[137]; 
    assign layer_0[273] = ~(in[149] ^ in[148]); 
    assign layer_0[274] = in[197] ^ in[195]; 
    assign layer_0[275] = in[91] | in[89]; 
    assign layer_0[276] = ~(in[136] | in[35]); 
    assign layer_0[277] = in[117] ^ in[155]; 
    assign layer_0[278] = in[143] | in[214]; 
    assign layer_0[279] = in[154] & in[138]; 
    assign layer_0[280] = in[134] ^ in[37]; 
    assign layer_0[281] = ~(in[44] ^ in[46]); 
    assign layer_0[282] = ~in[251]; 
    assign layer_0[283] = in[152] | in[82]; 
    assign layer_0[284] = in[35]; 
    assign layer_0[285] = in[88] & ~in[168]; 
    assign layer_0[286] = ~in[123]; 
    assign layer_0[287] = ~(in[214] | in[246]); 
    assign layer_0[288] = ~in[131]; 
    assign layer_0[289] = in[23] ^ in[93]; 
    assign layer_0[290] = ~(in[171] ^ in[164]); 
    assign layer_0[291] = in[154] & ~in[213]; 
    assign layer_0[292] = in[8] | in[219]; 
    assign layer_0[293] = ~(in[103] | in[145]); 
    assign layer_0[294] = ~(in[85] | in[177]); 
    assign layer_0[295] = ~(in[57] ^ in[171]); 
    assign layer_0[296] = in[38] ^ in[103]; 
    assign layer_0[297] = ~in[203]; 
    assign layer_0[298] = ~in[189] | (in[148] & in[189]); 
    assign layer_0[299] = in[183] | in[242]; 
    assign layer_0[300] = in[101] ^ in[99]; 
    assign layer_0[301] = ~in[182] | (in[162] & in[182]); 
    assign layer_0[302] = ~in[133] | (in[244] & in[133]); 
    assign layer_0[303] = in[89] & ~in[85]; 
    assign layer_0[304] = ~in[146] | (in[138] & in[146]); 
    assign layer_0[305] = ~(in[184] ^ in[77]); 
    assign layer_0[306] = in[215] & ~in[51]; 
    assign layer_0[307] = in[178] | in[205]; 
    assign layer_0[308] = ~(in[170] ^ in[126]); 
    assign layer_0[309] = ~in[170] | (in[170] & in[119]); 
    assign layer_0[310] = in[75] ^ in[89]; 
    assign layer_0[311] = in[247] ^ in[218]; 
    assign layer_0[312] = ~in[217]; 
    assign layer_0[313] = ~(in[247] ^ in[250]); 
    assign layer_0[314] = in[27] ^ in[210]; 
    assign layer_0[315] = ~in[98]; 
    assign layer_0[316] = ~in[58] | (in[152] & in[58]); 
    assign layer_0[317] = ~(in[252] ^ in[120]); 
    assign layer_0[318] = ~(in[26] | in[171]); 
    assign layer_0[319] = in[114] | in[93]; 
    assign layer_0[320] = in[211] ^ in[246]; 
    assign layer_0[321] = in[38] ^ in[68]; 
    assign layer_0[322] = in[98]; 
    assign layer_0[323] = ~(in[142] | in[162]); 
    assign layer_0[324] = in[235] & in[170]; 
    assign layer_0[325] = ~in[145] | (in[238] & in[145]); 
    assign layer_0[326] = in[220] ^ in[196]; 
    assign layer_0[327] = in[44] ^ in[74]; 
    assign layer_0[328] = in[120]; 
    assign layer_0[329] = ~(in[106] ^ in[108]); 
    assign layer_0[330] = ~in[137] | (in[137] & in[179]); 
    assign layer_0[331] = in[54] ^ in[81]; 
    assign layer_0[332] = in[163] & ~in[231]; 
    assign layer_0[333] = ~(in[183] ^ in[180]); 
    assign layer_0[334] = ~in[150]; 
    assign layer_0[335] = in[106] ^ in[58]; 
    assign layer_0[336] = ~(in[131] ^ in[121]); 
    assign layer_0[337] = in[146] ^ in[136]; 
    assign layer_0[338] = in[27] ^ in[87]; 
    assign layer_0[339] = in[165] | in[167]; 
    assign layer_0[340] = in[245] ^ in[214]; 
    assign layer_0[341] = ~(in[231] | in[248]); 
    assign layer_0[342] = in[57] & ~in[121]; 
    assign layer_0[343] = in[232]; 
    assign layer_0[344] = in[228] ^ in[197]; 
    assign layer_0[345] = ~(in[141] | in[142]); 
    assign layer_0[346] = in[99] ^ in[68]; 
    assign layer_0[347] = ~in[39] | (in[39] & in[148]); 
    assign layer_0[348] = ~in[183] | (in[183] & in[155]); 
    assign layer_0[349] = ~(in[20] | in[69]); 
    assign layer_0[350] = in[217] | in[61]; 
    assign layer_0[351] = in[131]; 
    assign layer_0[352] = in[71] ^ in[213]; 
    assign layer_0[353] = ~(in[241] | in[105]); 
    assign layer_0[354] = ~(in[56] ^ in[25]); 
    assign layer_0[355] = ~(in[199] ^ in[29]); 
    assign layer_0[356] = ~(in[228] ^ in[197]); 
    assign layer_0[357] = ~in[153] | (in[153] & in[204]); 
    assign layer_0[358] = in[197] & ~in[193]; 
    assign layer_0[359] = ~(in[99] | in[54]); 
    assign layer_0[360] = in[115] | in[83]; 
    assign layer_0[361] = ~(in[111] ^ in[109]); 
    assign layer_0[362] = ~(in[106] & in[56]); 
    assign layer_0[363] = in[95] ^ in[30]; 
    assign layer_0[364] = in[200]; 
    assign layer_0[365] = in[83] ^ in[52]; 
    assign layer_0[366] = ~in[153]; 
    assign layer_0[367] = ~in[24]; 
    assign layer_0[368] = ~(in[142] ^ in[45]); 
    assign layer_0[369] = in[44] | in[195]; 
    assign layer_0[370] = in[192] | in[219]; 
    assign layer_0[371] = in[197] | in[198]; 
    assign layer_0[372] = in[230] ^ in[183]; 
    assign layer_0[373] = in[124] ^ in[155]; 
    assign layer_0[374] = in[231] & ~in[179]; 
    assign layer_0[375] = ~(in[105] ^ in[194]); 
    assign layer_0[376] = ~(in[182] ^ in[155]); 
    assign layer_0[377] = ~(in[40] ^ in[89]); 
    assign layer_0[378] = ~(in[237] | in[147]); 
    assign layer_0[379] = in[76] ^ in[77]; 
    assign layer_0[380] = in[245] ^ in[113]; 
    assign layer_0[381] = ~(in[58] ^ in[249]); 
    assign layer_0[382] = ~(in[134] ^ in[164]); 
    assign layer_0[383] = ~(in[185] ^ in[67]); 
    assign layer_0[384] = ~(in[91] | in[66]); 
    assign layer_0[385] = ~(in[121] ^ in[154]); 
    assign layer_0[386] = in[119] ^ in[149]; 
    assign layer_0[387] = ~in[104] | (in[204] & in[104]); 
    assign layer_0[388] = ~(in[244] ^ in[198]); 
    assign layer_0[389] = ~(in[213] ^ in[228]); 
    assign layer_0[390] = ~(in[149] ^ in[147]); 
    assign layer_0[391] = in[215] ^ in[228]; 
    assign layer_0[392] = ~(in[218] | in[234]); 
    assign layer_0[393] = ~(in[182] ^ in[164]); 
    assign layer_0[394] = ~(in[22] | in[52]); 
    assign layer_0[395] = ~(in[131] | in[133]); 
    assign layer_0[396] = in[72] ^ in[28]; 
    assign layer_0[397] = in[27] ^ in[20]; 
    assign layer_0[398] = in[53]; 
    assign layer_0[399] = in[101]; 
    assign layer_0[400] = ~in[106]; 
    assign layer_0[401] = in[252] | in[183]; 
    assign layer_0[402] = in[220] ^ in[87]; 
    assign layer_0[403] = ~in[212] | (in[188] & in[212]); 
    assign layer_0[404] = in[118]; 
    assign layer_0[405] = ~(in[10] | in[86]); 
    assign layer_0[406] = ~(in[121] ^ in[171]); 
    assign layer_0[407] = in[41]; 
    assign layer_0[408] = in[148] | in[220]; 
    assign layer_0[409] = ~(in[89] ^ in[92]); 
    assign layer_0[410] = in[40] ^ in[98]; 
    assign layer_0[411] = ~(in[6] | in[177]); 
    assign layer_0[412] = ~in[135] | (in[135] & in[165]); 
    assign layer_0[413] = ~(in[131] | in[132]); 
    assign layer_0[414] = in[137] ^ in[10]; 
    assign layer_0[415] = ~in[211]; 
    assign layer_0[416] = ~in[100]; 
    assign layer_0[417] = in[101] ^ in[57]; 
    assign layer_0[418] = in[130] ^ in[163]; 
    assign layer_0[419] = ~(in[169] ^ in[157]); 
    assign layer_0[420] = in[137] | in[138]; 
    assign layer_0[421] = ~(in[196] ^ in[198]); 
    assign layer_0[422] = ~(in[9] | in[218]); 
    assign layer_0[423] = in[168] & ~in[95]; 
    assign layer_0[424] = ~(in[122] ^ in[155]); 
    assign layer_0[425] = in[219] ^ in[251]; 
    assign layer_0[426] = in[167] & ~in[177]; 
    assign layer_0[427] = in[237] | in[206]; 
    assign layer_0[428] = ~(in[59] ^ in[38]); 
    assign layer_0[429] = in[124] & ~in[199]; 
    assign layer_0[430] = in[167]; 
    assign layer_0[431] = ~(in[52] ^ in[58]); 
    assign layer_0[432] = ~(in[75] ^ in[106]); 
    assign layer_0[433] = in[229]; 
    assign layer_0[434] = ~(in[111] ^ in[109]); 
    assign layer_0[435] = in[53] & ~in[200]; 
    assign layer_0[436] = in[10] & ~in[75]; 
    assign layer_0[437] = ~(in[230] ^ in[248]); 
    assign layer_0[438] = ~(in[88] ^ in[58]); 
    assign layer_0[439] = ~(in[138] ^ in[172]); 
    assign layer_0[440] = in[93] | in[99]; 
    assign layer_0[441] = ~(in[72] ^ in[45]); 
    assign layer_0[442] = ~(in[100] ^ in[98]); 
    assign layer_0[443] = in[197] ^ in[166]; 
    assign layer_0[444] = ~(in[163] ^ in[133]); 
    assign layer_0[445] = ~(in[117] ^ in[103]); 
    assign layer_0[446] = in[146] ^ in[148]; 
    assign layer_0[447] = in[86] & ~in[181]; 
    assign layer_0[448] = in[116] ^ in[114]; 
    assign layer_0[449] = in[245] ^ in[196]; 
    assign layer_0[450] = in[153]; 
    assign layer_0[451] = ~(in[131] | in[76]); 
    assign layer_0[452] = ~in[38]; 
    assign layer_0[453] = ~(in[162] | in[163]); 
    assign layer_0[454] = in[169] & ~in[197]; 
    assign layer_0[455] = ~in[149] | (in[47] & in[149]); 
    assign layer_0[456] = in[59] ^ in[125]; 
    assign layer_0[457] = ~in[59] | (in[59] & in[122]); 
    assign layer_0[458] = in[108] ^ in[125]; 
    assign layer_0[459] = ~in[35]; 
    assign layer_0[460] = in[216] ^ in[68]; 
    assign layer_0[461] = ~(in[220] | in[27]); 
    assign layer_0[462] = in[124] | in[156]; 
    assign layer_0[463] = ~(in[100] | in[102]); 
    assign layer_0[464] = ~(in[195] | in[40]); 
    assign layer_0[465] = ~(in[250] | in[165]); 
    assign layer_0[466] = in[37] ^ in[51]; 
    assign layer_0[467] = in[155]; 
    assign layer_0[468] = ~in[26]; 
    assign layer_0[469] = ~(in[132] ^ in[146]); 
    assign layer_0[470] = in[201] | in[180]; 
    assign layer_0[471] = ~(in[237] ^ in[30]); 
    assign layer_0[472] = ~(in[189] ^ in[209]); 
    assign layer_0[473] = ~(in[194] | in[199]); 
    assign layer_0[474] = ~(in[203] | in[140]); 
    assign layer_0[475] = ~(in[165] ^ in[135]); 
    assign layer_0[476] = in[194] | in[26]; 
    assign layer_0[477] = ~(in[156] | in[122]); 
    assign layer_0[478] = ~(in[49] | in[92]); 
    assign layer_0[479] = in[21] ^ in[52]; 
    assign layer_0[480] = in[114] | in[165]; 
    assign layer_0[481] = in[213]; 
    assign layer_0[482] = ~(in[76] ^ in[120]); 
    assign layer_0[483] = ~in[198] | (in[198] & in[77]); 
    assign layer_0[484] = ~(in[86] ^ in[103]); 
    assign layer_0[485] = ~in[71] | (in[156] & in[71]); 
    assign layer_0[486] = ~(in[170] | in[139]); 
    assign layer_0[487] = in[88]; 
    assign layer_0[488] = in[21] ^ in[53]; 
    assign layer_0[489] = ~(in[83] ^ in[167]); 
    assign layer_0[490] = in[61] & in[108]; 
    assign layer_0[491] = in[197] ^ in[232]; 
    assign layer_0[492] = ~(in[108] | in[35]); 
    assign layer_0[493] = in[46] ^ in[169]; 
    assign layer_0[494] = in[55] ^ in[86]; 
    assign layer_0[495] = ~(in[216] ^ in[250]); 
    assign layer_0[496] = in[120] ^ in[166]; 
    assign layer_0[497] = ~(in[93] ^ in[63]); 
    assign layer_0[498] = ~(in[83] ^ in[202]); 
    assign layer_0[499] = in[84] ^ in[98]; 
    assign layer_0[500] = ~(in[101] | in[170]); 
    assign layer_0[501] = in[183] | in[147]; 
    assign layer_0[502] = ~(in[251] | in[186]); 
    assign layer_0[503] = in[40] & ~in[124]; 
    assign layer_0[504] = in[158] | in[215]; 
    assign layer_0[505] = ~(in[89] | in[72]); 
    assign layer_0[506] = ~in[143]; 
    assign layer_0[507] = in[118] & ~in[116]; 
    assign layer_0[508] = ~(in[214] ^ in[245]); 
    assign layer_0[509] = in[22] ^ in[214]; 
    assign layer_0[510] = in[70] ^ in[38]; 
    assign layer_0[511] = ~(in[97] | in[136]); 
    assign layer_0[512] = in[58] ^ in[29]; 
    assign layer_0[513] = in[91] & ~in[88]; 
    assign layer_0[514] = in[166] ^ in[244]; 
    assign layer_0[515] = in[63] | in[46]; 
    assign layer_0[516] = ~(in[216] ^ in[247]); 
    assign layer_0[517] = in[243] | in[12]; 
    assign layer_0[518] = ~(in[163] ^ in[158]); 
    assign layer_0[519] = in[120] & ~in[172]; 
    assign layer_0[520] = ~(in[37] ^ in[104]); 
    assign layer_0[521] = in[165] & ~in[26]; 
    assign layer_0[522] = ~(in[133] ^ in[147]); 
    assign layer_0[523] = ~(in[183] | in[158]); 
    assign layer_0[524] = ~(in[163] | in[165]); 
    assign layer_0[525] = ~(in[5] ^ in[6]); 
    assign layer_0[526] = in[56] & ~in[74]; 
    assign layer_0[527] = in[147] & ~in[231]; 
    assign layer_0[528] = in[151] & ~in[68]; 
    assign layer_0[529] = in[199] & ~in[164]; 
    assign layer_0[530] = in[19]; 
    assign layer_0[531] = ~(in[104] & in[152]); 
    assign layer_0[532] = in[114] | in[116]; 
    assign layer_0[533] = in[53] | in[38]; 
    assign layer_0[534] = ~(in[71] ^ in[59]); 
    assign layer_0[535] = in[246] ^ in[199]; 
    assign layer_0[536] = in[116] & in[107]; 
    assign layer_0[537] = ~in[171] | (in[171] & in[136]); 
    assign layer_0[538] = ~(in[101] ^ in[87]); 
    assign layer_0[539] = ~(in[242] | in[171]); 
    assign layer_0[540] = 1'b1; 
    assign layer_0[541] = ~(in[136] | in[245]); 
    assign layer_0[542] = in[222] ^ in[194]; 
    assign layer_0[543] = in[139] | in[178]; 
    assign layer_0[544] = ~(in[101] ^ in[113]); 
    assign layer_0[545] = ~(in[120] ^ in[50]); 
    assign layer_0[546] = in[45] ^ in[156]; 
    assign layer_0[547] = in[51] ^ in[246]; 
    assign layer_0[548] = ~(in[89] | in[58]); 
    assign layer_0[549] = in[136] & ~in[115]; 
    assign layer_0[550] = in[45]; 
    assign layer_0[551] = ~(in[59] ^ in[88]); 
    assign layer_0[552] = in[141]; 
    assign layer_0[553] = ~(in[163] ^ in[115]); 
    assign layer_0[554] = in[202]; 
    assign layer_0[555] = in[175] ^ in[178]; 
    assign layer_0[556] = ~(in[196] ^ in[38]); 
    assign layer_0[557] = ~(in[142] | in[165]); 
    assign layer_0[558] = in[89] ^ in[211]; 
    assign layer_0[559] = in[57] | in[88]; 
    assign layer_0[560] = in[131]; 
    assign layer_0[561] = ~(in[151] & in[166]); 
    assign layer_0[562] = ~(in[8] | in[28]); 
    assign layer_0[563] = in[115] & ~in[59]; 
    assign layer_0[564] = in[204] | in[192]; 
    assign layer_0[565] = in[155] ^ in[92]; 
    assign layer_0[566] = in[200] | in[28]; 
    assign layer_0[567] = ~(in[221] ^ in[152]); 
    assign layer_0[568] = in[155] | in[242]; 
    assign layer_0[569] = in[154] & ~in[179]; 
    assign layer_0[570] = ~in[85] | (in[147] & in[85]); 
    assign layer_0[571] = in[118] | in[112]; 
    assign layer_0[572] = in[20] ^ in[7]; 
    assign layer_0[573] = in[59] ^ in[235]; 
    assign layer_0[574] = in[201] | in[52]; 
    assign layer_0[575] = ~(in[11] | in[52]); 
    assign layer_0[576] = in[87] | in[132]; 
    assign layer_0[577] = ~(in[148] ^ in[146]); 
    assign layer_0[578] = ~in[46]; 
    assign layer_0[579] = ~in[100] | (in[171] & in[100]); 
    assign layer_0[580] = in[228] ^ in[233]; 
    assign layer_0[581] = ~(in[131] ^ in[178]); 
    assign layer_0[582] = ~(in[167] | in[237]); 
    assign layer_0[583] = in[186] ^ in[155]; 
    assign layer_0[584] = in[47] | in[177]; 
    assign layer_0[585] = ~(in[230] ^ in[44]); 
    assign layer_0[586] = in[29] ^ in[62]; 
    assign layer_0[587] = ~in[147] | (in[68] & in[147]); 
    assign layer_0[588] = in[147] ^ in[149]; 
    assign layer_0[589] = in[134] & ~in[147]; 
    assign layer_0[590] = ~(in[165] ^ in[136]); 
    assign layer_0[591] = in[129] | in[147]; 
    assign layer_0[592] = ~(in[151] | in[120]); 
    assign layer_0[593] = ~(in[141] | in[19]); 
    assign layer_0[594] = ~(in[72] ^ in[76]); 
    assign layer_0[595] = ~(in[92] ^ in[155]); 
    assign layer_0[596] = in[118]; 
    assign layer_0[597] = in[54] ^ in[105]; 
    assign layer_0[598] = in[39] & ~in[87]; 
    assign layer_0[599] = ~(in[185] ^ in[155]); 
    assign layer_0[600] = in[83] | in[52]; 
    assign layer_0[601] = ~(in[70] ^ in[201]); 
    assign layer_0[602] = ~(in[59] | in[75]); 
    assign layer_0[603] = ~(in[119] ^ in[90]); 
    assign layer_0[604] = ~(in[233] ^ in[202]); 
    assign layer_0[605] = in[250] | in[232]; 
    assign layer_0[606] = ~(in[150] | in[166]); 
    assign layer_0[607] = ~(in[143] | in[213]); 
    assign layer_0[608] = ~(in[40] ^ in[187]); 
    assign layer_0[609] = in[117] ^ in[115]; 
    assign layer_0[610] = ~(in[114] | in[57]); 
    assign layer_0[611] = in[201] | in[232]; 
    assign layer_0[612] = in[11] | in[12]; 
    assign layer_0[613] = in[26] ^ in[27]; 
    assign layer_0[614] = ~(in[251] | in[137]); 
    assign layer_0[615] = in[217] & ~in[120]; 
    assign layer_0[616] = ~(in[154] ^ in[106]); 
    assign layer_0[617] = in[59] | in[98]; 
    assign layer_0[618] = in[165] ^ in[163]; 
    assign layer_0[619] = ~in[131] | (in[131] & in[150]); 
    assign layer_0[620] = ~in[245] | (in[214] & in[245]); 
    assign layer_0[621] = in[76]; 
    assign layer_0[622] = in[23] | in[210]; 
    assign layer_0[623] = ~in[170] | (in[170] & in[180]); 
    assign layer_0[624] = ~in[214] | (in[88] & in[214]); 
    assign layer_0[625] = in[228]; 
    assign layer_0[626] = in[123]; 
    assign layer_0[627] = ~(in[121] | in[136]); 
    assign layer_0[628] = in[120]; 
    assign layer_0[629] = ~(in[61] ^ in[237]); 
    assign layer_0[630] = in[232] & in[105]; 
    assign layer_0[631] = in[161] | in[199]; 
    assign layer_0[632] = ~(in[243] ^ in[247]); 
    assign layer_0[633] = in[114]; 
    assign layer_0[634] = in[98] ^ in[83]; 
    assign layer_0[635] = in[41] ^ in[9]; 
    assign layer_0[636] = ~(in[230] ^ in[199]); 
    assign layer_0[637] = in[58] & ~in[27]; 
    assign layer_0[638] = ~(in[69] ^ in[151]); 
    assign layer_0[639] = ~in[153] | (in[153] & in[219]); 
    assign layer_0[640] = ~(in[110] ^ in[109]); 
    assign layer_0[641] = in[154] ^ in[172]; 
    assign layer_0[642] = in[233]; 
    assign layer_0[643] = ~in[136]; 
    assign layer_0[644] = in[163] & ~in[120]; 
    assign layer_0[645] = ~(in[177] | in[134]); 
    assign layer_0[646] = ~(in[178] ^ in[180]); 
    assign layer_0[647] = in[87] & ~in[44]; 
    assign layer_0[648] = in[151]; 
    assign layer_0[649] = in[158] | in[24]; 
    assign layer_0[650] = in[146] | in[139]; 
    assign layer_0[651] = in[164] ^ in[138]; 
    assign layer_0[652] = in[120] & ~in[101]; 
    assign layer_0[653] = ~in[215] | (in[138] & in[215]); 
    assign layer_0[654] = ~in[25] | (in[91] & in[25]); 
    assign layer_0[655] = in[135] ^ in[152]; 
    assign layer_0[656] = in[141] | in[123]; 
    assign layer_0[657] = in[236] ^ in[22]; 
    assign layer_0[658] = in[105] | in[28]; 
    assign layer_0[659] = in[107] | in[139]; 
    assign layer_0[660] = ~(in[98] ^ in[93]); 
    assign layer_0[661] = ~in[137]; 
    assign layer_0[662] = ~in[199] | (in[194] & in[199]); 
    assign layer_0[663] = in[104] | in[34]; 
    assign layer_0[664] = ~(in[103] ^ in[107]); 
    assign layer_0[665] = in[65] ^ in[19]; 
    assign layer_0[666] = ~(in[125] ^ in[105]); 
    assign layer_0[667] = 1'b0; 
    assign layer_0[668] = in[252]; 
    assign layer_0[669] = in[141] | in[214]; 
    assign layer_0[670] = in[59] ^ in[27]; 
    assign layer_0[671] = in[90]; 
    assign layer_0[672] = in[141] | in[250]; 
    assign layer_0[673] = ~(in[99] ^ in[113]); 
    assign layer_0[674] = ~(in[233] ^ in[231]); 
    assign layer_0[675] = ~(in[205] | in[203]); 
    assign layer_0[676] = ~(in[52] ^ in[200]); 
    assign layer_0[677] = ~in[248] | (in[248] & in[122]); 
    assign layer_0[678] = ~in[72] | (in[187] & in[72]); 
    assign layer_0[679] = in[26] | in[20]; 
    assign layer_0[680] = ~(in[129] ^ in[115]); 
    assign layer_0[681] = in[134] & ~in[136]; 
    assign layer_0[682] = in[199] ^ in[44]; 
    assign layer_0[683] = ~(in[163] | in[28]); 
    assign layer_0[684] = in[168] | in[23]; 
    assign layer_0[685] = ~(in[58] | in[194]); 
    assign layer_0[686] = ~(in[69] ^ in[89]); 
    assign layer_0[687] = in[104] | in[133]; 
    assign layer_0[688] = ~(in[173] | in[145]); 
    assign layer_0[689] = ~(in[186] ^ in[234]); 
    assign layer_0[690] = in[165] & ~in[127]; 
    assign layer_0[691] = in[141] | in[34]; 
    assign layer_0[692] = ~(in[31] ^ in[121]); 
    assign layer_0[693] = in[24] ^ in[72]; 
    assign layer_0[694] = ~(in[162] ^ in[215]); 
    assign layer_0[695] = ~in[105]; 
    assign layer_0[696] = in[138] ^ in[169]; 
    assign layer_0[697] = in[27] ^ in[72]; 
    assign layer_0[698] = ~(in[124] | in[83]); 
    assign layer_0[699] = in[180] | in[182]; 
    assign layer_0[700] = in[164] ^ in[135]; 
    assign layer_0[701] = in[210] ^ in[243]; 
    assign layer_0[702] = ~in[114]; 
    assign layer_0[703] = in[29] | in[104]; 
    assign layer_0[704] = ~(in[27] ^ in[73]); 
    assign layer_0[705] = in[158] ^ in[118]; 
    assign layer_0[706] = ~(in[162] ^ in[100]); 
    assign layer_0[707] = in[138] & ~in[106]; 
    assign layer_0[708] = in[214] ^ in[151]; 
    assign layer_0[709] = in[243] & ~in[231]; 
    assign layer_0[710] = in[211] ^ in[88]; 
    assign layer_0[711] = ~in[71]; 
    assign layer_0[712] = in[93] ^ in[91]; 
    assign layer_0[713] = ~(in[162] ^ in[164]); 
    assign layer_0[714] = in[40] ^ in[24]; 
    assign layer_0[715] = in[110] | in[78]; 
    assign layer_0[716] = ~(in[243] | in[101]); 
    assign layer_0[717] = ~(in[143] ^ in[242]); 
    assign layer_0[718] = ~in[73]; 
    assign layer_0[719] = in[203] | in[184]; 
    assign layer_0[720] = ~(in[234] ^ in[181]); 
    assign layer_0[721] = ~(in[91] ^ in[88]); 
    assign layer_0[722] = ~in[53]; 
    assign layer_0[723] = ~(in[105] | in[105]); 
    assign layer_0[724] = in[181] ^ in[164]; 
    assign layer_0[725] = ~in[74] | (in[74] & in[233]); 
    assign layer_0[726] = in[61] ^ in[44]; 
    assign layer_0[727] = ~(in[211] ^ in[196]); 
    assign layer_0[728] = ~(in[91] | in[92]); 
    assign layer_0[729] = ~in[162]; 
    assign layer_0[730] = in[137] & ~in[101]; 
    assign layer_0[731] = in[91] & ~in[26]; 
    assign layer_0[732] = ~(in[89] | in[171]); 
    assign layer_0[733] = in[250] ^ in[165]; 
    assign layer_0[734] = ~in[168]; 
    assign layer_0[735] = in[70]; 
    assign layer_0[736] = in[36] ^ in[79]; 
    assign layer_0[737] = ~(in[86] ^ in[74]); 
    assign layer_0[738] = in[47]; 
    assign layer_0[739] = ~(in[157] | in[140]); 
    assign layer_0[740] = in[38] & ~in[130]; 
    assign layer_0[741] = ~(in[87] ^ in[101]); 
    assign layer_0[742] = in[118] & ~in[219]; 
    assign layer_0[743] = ~(in[53] | in[83]); 
    assign layer_0[744] = ~(in[69] ^ in[67]); 
    assign layer_0[745] = in[235] & ~in[93]; 
    assign layer_0[746] = ~(in[140] | in[126]); 
    assign layer_0[747] = ~in[184] | (in[37] & in[184]); 
    assign layer_0[748] = ~(in[123] ^ in[141]); 
    assign layer_0[749] = in[219] & ~in[165]; 
    assign layer_0[750] = in[155] & in[139]; 
    assign layer_0[751] = in[85] & ~in[34]; 
    assign layer_0[752] = in[100] ^ in[200]; 
    assign layer_0[753] = ~(in[59] ^ in[87]); 
    assign layer_0[754] = ~(in[252] | in[245]); 
    assign layer_0[755] = ~(in[109] ^ in[106]); 
    assign layer_0[756] = ~(in[93] | in[111]); 
    assign layer_0[757] = in[52] | in[63]; 
    assign layer_0[758] = ~(in[197] | in[142]); 
    assign layer_0[759] = in[74] | in[61]; 
    assign layer_0[760] = ~(in[245] ^ in[198]); 
    assign layer_0[761] = ~(in[174] | in[9]); 
    assign layer_0[762] = ~in[127]; 
    assign layer_0[763] = ~(in[54] ^ in[99]); 
    assign layer_0[764] = in[46] ^ in[29]; 
    assign layer_0[765] = ~in[102] | (in[102] & in[24]); 
    assign layer_0[766] = ~(in[189] | in[219]); 
    assign layer_0[767] = ~(in[98] ^ in[81]); 
    assign layer_0[768] = ~(in[41] | in[192]); 
    assign layer_0[769] = in[106] & ~in[119]; 
    assign layer_0[770] = in[243] ^ in[211]; 
    assign layer_0[771] = in[206] ^ in[21]; 
    assign layer_0[772] = in[35] ^ in[21]; 
    assign layer_0[773] = in[134] ^ in[103]; 
    assign layer_0[774] = ~(in[13] ^ in[38]); 
    assign layer_0[775] = in[216] ^ in[103]; 
    assign layer_0[776] = in[116]; 
    assign layer_0[777] = ~(in[108] | in[26]); 
    assign layer_0[778] = in[73]; 
    assign layer_0[779] = in[92] & ~in[117]; 
    assign layer_0[780] = ~in[53]; 
    assign layer_0[781] = in[132] ^ in[102]; 
    assign layer_0[782] = in[83]; 
    assign layer_0[783] = ~(in[107] | in[139]); 
    assign layer_0[784] = ~(in[158] | in[111]); 
    assign layer_0[785] = in[120] & ~in[65]; 
    assign layer_0[786] = in[182] ^ in[196]; 
    assign layer_0[787] = in[172] | in[89]; 
    assign layer_0[788] = ~(in[151] ^ in[149]); 
    assign layer_0[789] = ~(in[168] ^ in[120]); 
    assign layer_0[790] = ~(in[195] ^ in[217]); 
    assign layer_0[791] = in[185] | in[232]; 
    assign layer_0[792] = ~(in[172] | in[251]); 
    assign layer_0[793] = in[72] ^ in[52]; 
    assign layer_0[794] = ~(in[157] ^ in[122]); 
    assign layer_0[795] = ~(in[182] | in[163]); 
    assign layer_0[796] = ~(in[119] ^ in[247]); 
    assign layer_0[797] = ~(in[170] ^ in[181]); 
    assign layer_0[798] = ~in[183] | (in[183] & in[91]); 
    assign layer_0[799] = in[61] ^ in[213]; 
    assign layer_0[800] = in[12]; 
    assign layer_0[801] = ~in[113] | (in[113] & in[205]); 
    assign layer_0[802] = in[102] & in[168]; 
    assign layer_0[803] = ~(in[234] ^ in[219]); 
    assign layer_0[804] = ~(in[119] | in[95]); 
    assign layer_0[805] = in[40] ^ in[42]; 
    assign layer_0[806] = ~(in[54] ^ in[74]); 
    assign layer_0[807] = in[40]; 
    assign layer_0[808] = in[103] & ~in[36]; 
    assign layer_0[809] = ~(in[251] | in[168]); 
    assign layer_0[810] = in[129] ^ in[243]; 
    assign layer_0[811] = ~(in[98] | in[105]); 
    assign layer_0[812] = in[114]; 
    assign layer_0[813] = ~(in[59] ^ in[57]); 
    assign layer_0[814] = ~(in[103] ^ in[132]); 
    assign layer_0[815] = ~(in[148] ^ in[165]); 
    assign layer_0[816] = ~in[215] | (in[183] & in[215]); 
    assign layer_0[817] = in[231] & ~in[164]; 
    assign layer_0[818] = in[40] & ~in[44]; 
    assign layer_0[819] = ~(in[8] | in[106]); 
    assign layer_0[820] = in[73] ^ in[97]; 
    assign layer_0[821] = ~(in[187] ^ in[196]); 
    assign layer_0[822] = ~in[93] | (in[93] & in[149]); 
    assign layer_0[823] = in[104] & ~in[72]; 
    assign layer_0[824] = ~(in[242] ^ in[203]); 
    assign layer_0[825] = ~(in[119] ^ in[90]); 
    assign layer_0[826] = in[92] | in[78]; 
    assign layer_0[827] = in[106] ^ in[94]; 
    assign layer_0[828] = ~(in[221] | in[41]); 
    assign layer_0[829] = ~in[133]; 
    assign layer_0[830] = in[47]; 
    assign layer_0[831] = in[152] ^ in[182]; 
    assign layer_0[832] = in[213] ^ in[23]; 
    assign layer_0[833] = ~in[201]; 
    assign layer_0[834] = ~in[151] | (in[151] & in[197]); 
    assign layer_0[835] = ~in[74] | (in[74] & in[72]); 
    assign layer_0[836] = in[9] & ~in[42]; 
    assign layer_0[837] = in[86] ^ in[221]; 
    assign layer_0[838] = in[52] | in[41]; 
    assign layer_0[839] = in[121] | in[137]; 
    assign layer_0[840] = in[136] | in[41]; 
    assign layer_0[841] = in[201] | in[248]; 
    assign layer_0[842] = ~(in[104] ^ in[251]); 
    assign layer_0[843] = ~(in[233] ^ in[105]); 
    assign layer_0[844] = ~(in[54] ^ in[58]); 
    assign layer_0[845] = ~(in[120] ^ in[83]); 
    assign layer_0[846] = ~(in[211] ^ in[197]); 
    assign layer_0[847] = in[180] ^ in[150]; 
    assign layer_0[848] = ~(in[61] ^ in[27]); 
    assign layer_0[849] = ~in[102] | (in[197] & in[102]); 
    assign layer_0[850] = in[101]; 
    assign layer_0[851] = ~(in[137] | in[247]); 
    assign layer_0[852] = ~(in[100] ^ in[86]); 
    assign layer_0[853] = in[138] & ~in[180]; 
    assign layer_0[854] = ~(in[57] ^ in[59]); 
    assign layer_0[855] = in[219]; 
    assign layer_0[856] = ~in[121] | (in[146] & in[121]); 
    assign layer_0[857] = in[213] ^ in[182]; 
    assign layer_0[858] = in[118] | in[232]; 
    assign layer_0[859] = ~(in[138] | in[19]); 
    assign layer_0[860] = in[221] ^ in[170]; 
    assign layer_0[861] = in[5] | in[172]; 
    assign layer_0[862] = in[103] ^ in[54]; 
    assign layer_0[863] = in[120] & ~in[148]; 
    assign layer_0[864] = in[183] | in[147]; 
    assign layer_0[865] = in[221] | in[228]; 
    assign layer_0[866] = ~(in[52] ^ in[81]); 
    assign layer_0[867] = in[243] | in[21]; 
    assign layer_0[868] = in[135] & ~in[86]; 
    assign layer_0[869] = in[8] & ~in[155]; 
    assign layer_0[870] = in[26] ^ in[60]; 
    assign layer_0[871] = in[75] | in[73]; 
    assign layer_0[872] = in[65] ^ in[83]; 
    assign layer_0[873] = ~(in[107] ^ in[87]); 
    assign layer_0[874] = in[55] & ~in[60]; 
    assign layer_0[875] = ~(in[76] ^ in[74]); 
    assign layer_0[876] = in[198] & ~in[231]; 
    assign layer_0[877] = ~in[72] | (in[60] & in[72]); 
    assign layer_0[878] = ~in[179] | (in[134] & in[179]); 
    assign layer_0[879] = in[226] ^ in[33]; 
    assign layer_0[880] = in[246]; 
    assign layer_0[881] = ~(in[189] ^ in[102]); 
    assign layer_0[882] = ~(in[234] ^ in[203]); 
    assign layer_0[883] = in[77] & ~in[46]; 
    assign layer_0[884] = ~(in[156] | in[117]); 
    assign layer_0[885] = ~(in[219] | in[203]); 
    assign layer_0[886] = ~(in[92] | in[54]); 
    assign layer_0[887] = in[104]; 
    assign layer_0[888] = ~(in[162] ^ in[181]); 
    assign layer_0[889] = ~(in[138] ^ in[89]); 
    assign layer_0[890] = ~(in[121] ^ in[153]); 
    assign layer_0[891] = ~(in[120] | in[105]); 
    assign layer_0[892] = ~(in[130] | in[85]); 
    assign layer_0[893] = ~in[24] | (in[69] & in[24]); 
    assign layer_0[894] = in[119] & ~in[109]; 
    assign layer_0[895] = in[24]; 
    assign layer_0[896] = ~in[122] | (in[216] & in[122]); 
    assign layer_0[897] = ~(in[74] ^ in[31]); 
    assign layer_0[898] = in[183] ^ in[121]; 
    assign layer_0[899] = in[19] | in[105]; 
    assign layer_0[900] = in[42] ^ in[53]; 
    assign layer_0[901] = ~(in[166] ^ in[197]); 
    assign layer_0[902] = ~in[187] | (in[187] & in[154]); 
    assign layer_0[903] = in[65] | in[34]; 
    assign layer_0[904] = ~(in[30] ^ in[59]); 
    assign layer_0[905] = ~(in[165] | in[104]); 
    assign layer_0[906] = in[227] | in[247]; 
    assign layer_0[907] = in[101] | in[115]; 
    assign layer_0[908] = in[126] | in[11]; 
    assign layer_0[909] = ~in[120]; 
    assign layer_0[910] = ~(in[40] ^ in[166]); 
    assign layer_0[911] = ~(in[179] ^ in[198]); 
    assign layer_0[912] = in[73] ^ in[61]; 
    assign layer_0[913] = ~(in[156] ^ in[137]); 
    assign layer_0[914] = in[94] | in[66]; 
    assign layer_0[915] = in[147]; 
    assign layer_0[916] = ~(in[30] ^ in[63]); 
    assign layer_0[917] = in[108] ^ in[90]; 
    assign layer_0[918] = ~(in[156] ^ in[120]); 
    assign layer_0[919] = ~(in[140] ^ in[155]); 
    assign layer_0[920] = ~(in[193] | in[227]); 
    assign layer_0[921] = ~(in[35] ^ in[66]); 
    assign layer_0[922] = in[9] ^ in[27]; 
    assign layer_0[923] = ~in[119]; 
    assign layer_0[924] = in[102] ^ in[113]; 
    assign layer_0[925] = in[145] | in[179]; 
    assign layer_0[926] = in[151] ^ in[120]; 
    assign layer_0[927] = in[141] | in[156]; 
    assign layer_0[928] = ~in[150] | (in[150] & in[107]); 
    assign layer_0[929] = ~(in[187] ^ in[156]); 
    assign layer_0[930] = ~(in[28] ^ in[25]); 
    assign layer_0[931] = ~(in[181] ^ in[83]); 
    assign layer_0[932] = ~(in[78] ^ in[243]); 
    assign layer_0[933] = in[157] ^ in[214]; 
    assign layer_0[934] = ~(in[221] ^ in[212]); 
    assign layer_0[935] = in[27] ^ in[10]; 
    assign layer_0[936] = in[37] | in[229]; 
    assign layer_0[937] = in[104] & in[199]; 
    assign layer_0[938] = ~(in[152] | in[21]); 
    assign layer_0[939] = in[171] & ~in[205]; 
    assign layer_0[940] = in[54] & ~in[101]; 
    assign layer_0[941] = in[195] ^ in[10]; 
    assign layer_0[942] = in[147] ^ in[149]; 
    assign layer_0[943] = in[27] ^ in[60]; 
    assign layer_0[944] = ~in[58] | (in[156] & in[58]); 
    assign layer_0[945] = ~in[41] | (in[116] & in[41]); 
    assign layer_0[946] = ~in[184] | (in[213] & in[184]); 
    assign layer_0[947] = in[232] & ~in[54]; 
    assign layer_0[948] = in[186] ^ in[34]; 
    assign layer_0[949] = ~(in[152] | in[232]); 
    assign layer_0[950] = in[137] & ~in[20]; 
    assign layer_0[951] = ~(in[85] | in[141]); 
    assign layer_0[952] = ~in[41]; 
    assign layer_0[953] = in[82] | in[98]; 
    assign layer_0[954] = in[198] | in[179]; 
    assign layer_0[955] = ~(in[122] | in[156]); 
    assign layer_0[956] = in[22] ^ in[89]; 
    assign layer_0[957] = in[52] ^ in[82]; 
    assign layer_0[958] = in[73] & ~in[181]; 
    assign layer_0[959] = in[106] & ~in[93]; 
    assign layer_0[960] = in[12] ^ in[241]; 
    assign layer_0[961] = ~(in[59] ^ in[89]); 
    assign layer_0[962] = in[199] ^ in[186]; 
    assign layer_0[963] = in[57] | in[114]; 
    assign layer_0[964] = ~(in[129] | in[130]); 
    assign layer_0[965] = in[154] | in[182]; 
    assign layer_0[966] = ~(in[103] ^ in[242]); 
    assign layer_0[967] = in[116] ^ in[149]; 
    assign layer_0[968] = in[204] ^ in[25]; 
    assign layer_0[969] = ~(in[39] | in[92]); 
    assign layer_0[970] = ~(in[111] ^ in[28]); 
    assign layer_0[971] = in[40] & ~in[243]; 
    assign layer_0[972] = ~in[89] | (in[89] & in[76]); 
    assign layer_0[973] = ~in[152] | (in[152] & in[164]); 
    assign layer_0[974] = in[109] | in[136]; 
    assign layer_0[975] = in[108]; 
    assign layer_0[976] = in[250] | in[136]; 
    assign layer_0[977] = ~(in[104] ^ in[62]); 
    assign layer_0[978] = in[183]; 
    assign layer_0[979] = in[246]; 
    assign layer_0[980] = ~(in[206] ^ in[143]); 
    assign layer_0[981] = ~(in[156] | in[105]); 
    assign layer_0[982] = in[36] & ~in[68]; 
    assign layer_0[983] = ~(in[237] ^ in[196]); 
    assign layer_0[984] = in[79] | in[228]; 
    assign layer_0[985] = in[69] | in[67]; 
    assign layer_0[986] = ~in[138]; 
    assign layer_0[987] = in[171] | in[188]; 
    assign layer_0[988] = ~(in[54] | in[38]); 
    assign layer_0[989] = in[165] | in[178]; 
    assign layer_0[990] = in[244] ^ in[105]; 
    assign layer_0[991] = in[132] ^ in[146]; 
    assign layer_0[992] = in[252] ^ in[247]; 
    assign layer_0[993] = ~(in[88] ^ in[103]); 
    assign layer_0[994] = in[118] ^ in[141]; 
    assign layer_0[995] = in[154] | in[98]; 
    assign layer_0[996] = in[136] | in[131]; 
    assign layer_0[997] = ~(in[135] | in[210]); 
    assign layer_0[998] = in[244] ^ in[252]; 
    assign layer_0[999] = in[165] ^ in[196]; 
    assign layer_0[1000] = ~(in[5] | in[120]); 
    assign layer_0[1001] = ~(in[158] | in[214]); 
    assign layer_0[1002] = in[141] ^ in[232]; 
    assign layer_0[1003] = in[152] & ~in[37]; 
    assign layer_0[1004] = ~in[197] | (in[197] & in[154]); 
    assign layer_0[1005] = ~(in[89] | in[90]); 
    assign layer_0[1006] = in[74] ^ in[77]; 
    assign layer_0[1007] = ~in[114]; 
    assign layer_0[1008] = ~(in[45] ^ in[107]); 
    assign layer_0[1009] = ~(in[11] | in[207]); 
    assign layer_0[1010] = in[190] ^ in[79]; 
    assign layer_0[1011] = in[88] | in[228]; 
    assign layer_0[1012] = ~in[91] | (in[25] & in[91]); 
    assign layer_0[1013] = ~(in[179] | in[243]); 
    assign layer_0[1014] = ~(in[113] | in[185]); 
    assign layer_0[1015] = in[23] ^ in[70]; 
    assign layer_0[1016] = in[150] | in[148]; 
    assign layer_0[1017] = in[216] ^ in[51]; 
    assign layer_0[1018] = ~in[182] | (in[182] & in[90]); 
    assign layer_0[1019] = in[90] ^ in[86]; 
    assign layer_0[1020] = ~in[218] | (in[218] & in[90]); 
    assign layer_0[1021] = in[130] ^ in[131]; 
    assign layer_0[1022] = ~(in[92] ^ in[61]); 
    assign layer_0[1023] = ~(in[187] ^ in[209]); 
    assign layer_0[1024] = ~in[106] | (in[106] & in[89]); 
    assign layer_0[1025] = ~(in[102] ^ in[91]); 
    assign layer_0[1026] = in[215]; 
    assign layer_0[1027] = in[38]; 
    assign layer_0[1028] = ~in[215]; 
    assign layer_0[1029] = ~in[182]; 
    assign layer_0[1030] = in[104] | in[42]; 
    assign layer_0[1031] = in[8] & ~in[165]; 
    assign layer_0[1032] = in[169] & ~in[89]; 
    assign layer_0[1033] = ~(in[62] ^ in[74]); 
    assign layer_0[1034] = ~(in[104] ^ in[57]); 
    assign layer_0[1035] = ~(in[164] | in[147]); 
    assign layer_0[1036] = ~(in[196] | in[248]); 
    assign layer_0[1037] = in[250] | in[242]; 
    assign layer_0[1038] = ~in[132] | (in[228] & in[132]); 
    assign layer_0[1039] = in[73] ^ in[106]; 
    assign layer_0[1040] = ~(in[147] | in[173]); 
    assign layer_0[1041] = ~(in[236] ^ in[21]); 
    assign layer_0[1042] = ~(in[85] ^ in[21]); 
    assign layer_0[1043] = in[108] ^ in[110]; 
    assign layer_0[1044] = in[186] ^ in[166]; 
    assign layer_0[1045] = in[216] & ~in[210]; 
    assign layer_0[1046] = in[115] ^ in[87]; 
    assign layer_0[1047] = in[117] ^ in[122]; 
    assign layer_0[1048] = ~(in[165] ^ in[167]); 
    assign layer_0[1049] = in[140] ^ in[215]; 
    assign layer_0[1050] = in[151] & ~in[101]; 
    assign layer_0[1051] = in[50] | in[36]; 
    assign layer_0[1052] = ~(in[153] ^ in[122]); 
    assign layer_0[1053] = ~in[154] | (in[154] & in[53]); 
    assign layer_0[1054] = ~(in[186] ^ in[218]); 
    assign layer_0[1055] = in[153] & ~in[235]; 
    assign layer_0[1056] = in[105]; 
    assign layer_0[1057] = ~(in[129] | in[168]); 
    assign layer_0[1058] = ~(in[167] | in[207]); 
    assign layer_0[1059] = ~(in[150] | in[119]); 
    assign layer_0[1060] = ~in[85] | (in[119] & in[85]); 
    assign layer_0[1061] = ~in[87] | (in[104] & in[87]); 
    assign layer_0[1062] = in[73]; 
    assign layer_0[1063] = in[40] & ~in[47]; 
    assign layer_0[1064] = in[234]; 
    assign layer_0[1065] = ~in[217] | (in[217] & in[249]); 
    assign layer_0[1066] = in[203] & ~in[157]; 
    assign layer_0[1067] = in[253] | in[245]; 
    assign layer_0[1068] = in[183] ^ in[21]; 
    assign layer_0[1069] = ~(in[106] | in[138]); 
    assign layer_0[1070] = in[155] & ~in[204]; 
    assign layer_0[1071] = in[26] ^ in[27]; 
    assign layer_0[1072] = in[77] ^ in[60]; 
    assign layer_0[1073] = ~in[87]; 
    assign layer_0[1074] = in[204] ^ in[237]; 
    assign layer_0[1075] = ~(in[132] | in[131]); 
    assign layer_0[1076] = in[111] | in[230]; 
    assign layer_0[1077] = ~in[38] | (in[38] & in[88]); 
    assign layer_0[1078] = in[184] & ~in[228]; 
    assign layer_0[1079] = ~(in[198] ^ in[188]); 
    assign layer_0[1080] = ~(in[163] ^ in[63]); 
    assign layer_0[1081] = in[151] | in[176]; 
    assign layer_0[1082] = in[198] | in[185]; 
    assign layer_0[1083] = ~(in[27] ^ in[106]); 
    assign layer_0[1084] = in[76] | in[107]; 
    assign layer_0[1085] = ~in[60] | (in[194] & in[60]); 
    assign layer_0[1086] = in[101] | in[229]; 
    assign layer_0[1087] = ~in[72]; 
    assign layer_0[1088] = ~(in[52] | in[26]); 
    assign layer_0[1089] = in[117] & ~in[236]; 
    assign layer_0[1090] = in[98]; 
    assign layer_0[1091] = in[156] ^ in[209]; 
    assign layer_0[1092] = in[97] & ~in[99]; 
    assign layer_0[1093] = in[79] | in[73]; 
    assign layer_0[1094] = in[46] | in[236]; 
    assign layer_0[1095] = in[104] & ~in[76]; 
    assign layer_0[1096] = in[117] & ~in[94]; 
    assign layer_0[1097] = ~(in[92] ^ in[110]); 
    assign layer_0[1098] = ~(in[164] ^ in[168]); 
    assign layer_0[1099] = in[206]; 
    assign layer_0[1100] = ~(in[180] ^ in[204]); 
    assign layer_0[1101] = in[115]; 
    assign layer_0[1102] = in[57] & ~in[23]; 
    assign layer_0[1103] = in[102] ^ in[97]; 
    assign layer_0[1104] = ~(in[151] ^ in[182]); 
    assign layer_0[1105] = in[148]; 
    assign layer_0[1106] = ~(in[146] | in[101]); 
    assign layer_0[1107] = in[71] ^ in[85]; 
    assign layer_0[1108] = in[110] ^ in[108]; 
    assign layer_0[1109] = ~(in[72] | in[252]); 
    assign layer_0[1110] = ~(in[124] ^ in[155]); 
    assign layer_0[1111] = in[41] ^ in[117]; 
    assign layer_0[1112] = ~in[108] | (in[108] & in[143]); 
    assign layer_0[1113] = ~(in[58] ^ in[172]); 
    assign layer_0[1114] = ~in[66] | (in[42] & in[66]); 
    assign layer_0[1115] = in[223] | in[20]; 
    assign layer_0[1116] = ~in[125] | (in[218] & in[125]); 
    assign layer_0[1117] = in[77] | in[101]; 
    assign layer_0[1118] = ~in[93]; 
    assign layer_0[1119] = in[136] ^ in[206]; 
    assign layer_0[1120] = ~(in[88] | in[195]); 
    assign layer_0[1121] = ~(in[219] | in[249]); 
    assign layer_0[1122] = ~(in[219] ^ in[165]); 
    assign layer_0[1123] = ~in[201]; 
    assign layer_0[1124] = ~(in[126] ^ in[21]); 
    assign layer_0[1125] = in[251] | in[103]; 
    assign layer_0[1126] = ~(in[29] ^ in[11]); 
    assign layer_0[1127] = in[43] | in[27]; 
    assign layer_0[1128] = ~(in[150] | in[212]); 
    assign layer_0[1129] = in[166]; 
    assign layer_0[1130] = in[177]; 
    assign layer_0[1131] = in[52] | in[69]; 
    assign layer_0[1132] = ~(in[213] | in[116]); 
    assign layer_0[1133] = ~in[75] | (in[75] & in[84]); 
    assign layer_0[1134] = in[26] ^ in[28]; 
    assign layer_0[1135] = in[164] ^ in[166]; 
    assign layer_0[1136] = ~(in[54] | in[69]); 
    assign layer_0[1137] = ~in[169] | (in[26] & in[169]); 
    assign layer_0[1138] = ~(in[148] | in[20]); 
    assign layer_0[1139] = in[141] ^ in[127]; 
    assign layer_0[1140] = ~(in[19] ^ in[70]); 
    assign layer_0[1141] = in[250] ^ in[168]; 
    assign layer_0[1142] = in[39] | in[228]; 
    assign layer_0[1143] = ~in[153] | (in[153] & in[196]); 
    assign layer_0[1144] = in[181] & ~in[36]; 
    assign layer_0[1145] = in[148] | in[146]; 
    assign layer_0[1146] = in[42] ^ in[167]; 
    assign layer_0[1147] = ~(in[137] | in[176]); 
    assign layer_0[1148] = in[65]; 
    assign layer_0[1149] = in[194] | in[27]; 
    assign layer_0[1150] = ~(in[10] ^ in[132]); 
    assign layer_0[1151] = in[57] ^ in[71]; 
    assign layer_0[1152] = in[201]; 
    assign layer_0[1153] = in[107] ^ in[74]; 
    assign layer_0[1154] = in[139] & ~in[195]; 
    assign layer_0[1155] = ~(in[162] ^ in[62]); 
    assign layer_0[1156] = in[41]; 
    assign layer_0[1157] = ~(in[220] ^ in[189]); 
    assign layer_0[1158] = in[154] ^ in[90]; 
    assign layer_0[1159] = in[86]; 
    assign layer_0[1160] = in[103] | in[148]; 
    assign layer_0[1161] = ~(in[171] | in[158]); 
    assign layer_0[1162] = in[83] ^ in[86]; 
    assign layer_0[1163] = in[136] | in[136]; 
    assign layer_0[1164] = ~(in[182] ^ in[228]); 
    assign layer_0[1165] = in[58] | in[76]; 
    assign layer_0[1166] = in[90] ^ in[92]; 
    assign layer_0[1167] = in[180] ^ in[101]; 
    assign layer_0[1168] = ~(in[57] ^ in[130]); 
    assign layer_0[1169] = ~in[114]; 
    assign layer_0[1170] = ~in[98] | (in[229] & in[98]); 
    assign layer_0[1171] = in[205] | in[188]; 
    assign layer_0[1172] = ~in[100]; 
    assign layer_0[1173] = in[79] | in[98]; 
    assign layer_0[1174] = ~(in[76] ^ in[83]); 
    assign layer_0[1175] = in[138] ^ in[129]; 
    assign layer_0[1176] = ~(in[202] ^ in[251]); 
    assign layer_0[1177] = ~(in[229] ^ in[221]); 
    assign layer_0[1178] = in[28] ^ in[61]; 
    assign layer_0[1179] = ~(in[243] | in[186]); 
    assign layer_0[1180] = in[72] ^ in[105]; 
    assign layer_0[1181] = ~(in[23] | in[154]); 
    assign layer_0[1182] = ~(in[57] | in[62]); 
    assign layer_0[1183] = ~(in[94] ^ in[92]); 
    assign layer_0[1184] = ~(in[58] ^ in[45]); 
    assign layer_0[1185] = ~(in[173] ^ in[118]); 
    assign layer_0[1186] = ~(in[9] ^ in[27]); 
    assign layer_0[1187] = ~(in[198] | in[165]); 
    assign layer_0[1188] = in[88] ^ in[41]; 
    assign layer_0[1189] = in[125] | in[94]; 
    assign layer_0[1190] = in[148] & ~in[199]; 
    assign layer_0[1191] = in[103] & ~in[83]; 
    assign layer_0[1192] = in[123] ^ in[165]; 
    assign layer_0[1193] = in[167] & ~in[92]; 
    assign layer_0[1194] = ~in[203] | (in[203] & in[98]); 
    assign layer_0[1195] = ~(in[50] | in[242]); 
    assign layer_0[1196] = ~(in[24] | in[157]); 
    assign layer_0[1197] = in[115]; 
    assign layer_0[1198] = in[212] | in[95]; 
    assign layer_0[1199] = in[104] & ~in[173]; 
    assign layer_0[1200] = in[63] ^ in[99]; 
    assign layer_0[1201] = in[40] ^ in[75]; 
    assign layer_0[1202] = in[71] ^ in[41]; 
    assign layer_0[1203] = in[151]; 
    assign layer_0[1204] = ~(in[155] | in[36]); 
    assign layer_0[1205] = in[163] | in[87]; 
    assign layer_0[1206] = in[129] | in[154]; 
    assign layer_0[1207] = in[140]; 
    assign layer_0[1208] = ~(in[30] | in[185]); 
    assign layer_0[1209] = in[156] & ~in[85]; 
    assign layer_0[1210] = in[52] | in[91]; 
    assign layer_0[1211] = in[149] & ~in[137]; 
    assign layer_0[1212] = ~(in[91] ^ in[88]); 
    assign layer_0[1213] = in[203] ^ in[232]; 
    assign layer_0[1214] = in[132]; 
    assign layer_0[1215] = in[135] & ~in[43]; 
    assign layer_0[1216] = ~(in[22] | in[36]); 
    assign layer_0[1217] = ~in[24] | (in[123] & in[24]); 
    assign layer_0[1218] = in[142] ^ in[140]; 
    assign layer_0[1219] = ~in[88]; 
    assign layer_0[1220] = ~in[232] | (in[70] & in[232]); 
    assign layer_0[1221] = ~(in[107] | in[124]); 
    assign layer_0[1222] = ~(in[109] ^ in[91]); 
    assign layer_0[1223] = in[93]; 
    assign layer_0[1224] = in[212] | in[237]; 
    assign layer_0[1225] = in[187] & ~in[90]; 
    assign layer_0[1226] = ~(in[147] ^ in[165]); 
    assign layer_0[1227] = in[166] ^ in[100]; 
    assign layer_0[1228] = ~(in[236] | in[149]); 
    assign layer_0[1229] = in[38] | in[54]; 
    assign layer_0[1230] = in[131] | in[122]; 
    assign layer_0[1231] = ~(in[140] ^ in[104]); 
    assign layer_0[1232] = in[40] | in[56]; 
    assign layer_0[1233] = in[173] | in[117]; 
    assign layer_0[1234] = in[9] ^ in[245]; 
    assign layer_0[1235] = in[119] & ~in[86]; 
    assign layer_0[1236] = ~(in[242] | in[87]); 
    assign layer_0[1237] = ~(in[139] ^ in[107]); 
    assign layer_0[1238] = in[134] & ~in[53]; 
    assign layer_0[1239] = in[76] ^ in[21]; 
    assign layer_0[1240] = in[198]; 
    assign layer_0[1241] = ~(in[235] | in[147]); 
    assign layer_0[1242] = ~(in[42] ^ in[89]); 
    assign layer_0[1243] = ~(in[69] ^ in[38]); 
    assign layer_0[1244] = ~(in[150] | in[135]); 
    assign layer_0[1245] = ~(in[125] ^ in[205]); 
    assign layer_0[1246] = in[131]; 
    assign layer_0[1247] = in[90] ^ in[54]; 
    assign layer_0[1248] = in[166] ^ in[186]; 
    assign layer_0[1249] = in[76] & ~in[27]; 
    assign layer_0[1250] = in[46] | in[63]; 
    assign layer_0[1251] = ~(in[210] | in[72]); 
    assign layer_0[1252] = ~(in[78] ^ in[76]); 
    assign layer_0[1253] = in[166] ^ in[244]; 
    assign layer_0[1254] = ~(in[162] ^ in[120]); 
    assign layer_0[1255] = in[246]; 
    assign layer_0[1256] = ~(in[77] ^ in[73]); 
    assign layer_0[1257] = ~in[203] | (in[203] & in[81]); 
    assign layer_0[1258] = in[150] ^ in[148]; 
    assign layer_0[1259] = ~(in[137] | in[9]); 
    assign layer_0[1260] = in[9] ^ in[40]; 
    assign layer_0[1261] = in[25] ^ in[20]; 
    assign layer_0[1262] = ~(in[101] ^ in[115]); 
    assign layer_0[1263] = ~(in[70] ^ in[162]); 
    assign layer_0[1264] = ~(in[22] | in[50]); 
    assign layer_0[1265] = in[158] ^ in[251]; 
    assign layer_0[1266] = ~in[186]; 
    assign layer_0[1267] = ~(in[232] | in[201]); 
    assign layer_0[1268] = ~(in[143] ^ in[177]); 
    assign layer_0[1269] = in[88] ^ in[131]; 
    assign layer_0[1270] = in[190] ^ in[188]; 
    assign layer_0[1271] = in[95] ^ in[93]; 
    assign layer_0[1272] = ~in[153]; 
    assign layer_0[1273] = ~(in[21] ^ in[197]); 
    assign layer_0[1274] = in[131] ^ in[119]; 
    assign layer_0[1275] = in[83] ^ in[79]; 
    assign layer_0[1276] = in[30] | in[63]; 
    assign layer_0[1277] = in[92] ^ in[78]; 
    assign layer_0[1278] = ~in[109]; 
    assign layer_0[1279] = ~in[154] | (in[154] & in[210]); 
    assign layer_0[1280] = ~in[186]; 
    assign layer_0[1281] = ~in[12]; 
    assign layer_0[1282] = ~(in[90] ^ in[155]); 
    assign layer_0[1283] = ~(in[35] ^ in[200]); 
    assign layer_0[1284] = ~(in[115] | in[93]); 
    assign layer_0[1285] = ~(in[140] ^ in[105]); 
    assign layer_0[1286] = ~(in[30] ^ in[63]); 
    assign layer_0[1287] = ~(in[123] | in[183]); 
    assign layer_0[1288] = in[215] & ~in[6]; 
    assign layer_0[1289] = in[118] ^ in[132]; 
    assign layer_0[1290] = ~(in[77] ^ in[56]); 
    assign layer_0[1291] = in[215] ^ in[249]; 
    assign layer_0[1292] = ~(in[90] ^ in[126]); 
    assign layer_0[1293] = in[41] ^ in[73]; 
    assign layer_0[1294] = ~in[89] | (in[60] & in[89]); 
    assign layer_0[1295] = in[25] ^ in[22]; 
    assign layer_0[1296] = in[120] ^ in[136]; 
    assign layer_0[1297] = in[86] ^ in[100]; 
    assign layer_0[1298] = in[217] ^ in[218]; 
    assign layer_0[1299] = ~(in[92] ^ in[55]); 
    assign layer_0[1300] = ~in[168]; 
    assign layer_0[1301] = in[11] | in[46]; 
    assign layer_0[1302] = in[19]; 
    assign layer_0[1303] = ~(in[119] ^ in[97]); 
    assign layer_0[1304] = in[214] | in[126]; 
    assign layer_0[1305] = ~in[120]; 
    assign layer_0[1306] = ~(in[169] | in[159]); 
    assign layer_0[1307] = ~in[218] | (in[218] & in[147]); 
    assign layer_0[1308] = ~(in[125] ^ in[169]); 
    assign layer_0[1309] = ~(in[54] | in[172]); 
    assign layer_0[1310] = ~(in[198] ^ in[212]); 
    assign layer_0[1311] = ~(in[183] ^ in[218]); 
    assign layer_0[1312] = in[207] ^ in[150]; 
    assign layer_0[1313] = ~(in[10] | in[29]); 
    assign layer_0[1314] = in[101] | in[30]; 
    assign layer_0[1315] = ~(in[63] | in[68]); 
    assign layer_0[1316] = ~in[54] | (in[179] & in[54]); 
    assign layer_0[1317] = ~(in[90] ^ in[87]); 
    assign layer_0[1318] = in[102] | in[116]; 
    assign layer_0[1319] = ~(in[154] ^ in[166]); 
    assign layer_0[1320] = ~(in[203] | in[202]); 
    assign layer_0[1321] = ~(in[125] | in[123]); 
    assign layer_0[1322] = in[99] | in[139]; 
    assign layer_0[1323] = ~(in[102] ^ in[53]); 
    assign layer_0[1324] = ~(in[179] ^ in[181]); 
    assign layer_0[1325] = in[67] ^ in[19]; 
    assign layer_0[1326] = in[230] ^ in[165]; 
    assign layer_0[1327] = ~(in[148] ^ in[119]); 
    assign layer_0[1328] = in[212]; 
    assign layer_0[1329] = in[163] | in[131]; 
    assign layer_0[1330] = ~(in[201] ^ in[198]); 
    assign layer_0[1331] = in[226] ^ in[196]; 
    assign layer_0[1332] = ~in[169]; 
    assign layer_0[1333] = ~(in[212] ^ in[77]); 
    assign layer_0[1334] = in[45] ^ in[78]; 
    assign layer_0[1335] = ~(in[51] ^ in[22]); 
    assign layer_0[1336] = in[19]; 
    assign layer_0[1337] = ~(in[114] | in[113]); 
    assign layer_0[1338] = in[67] ^ in[35]; 
    assign layer_0[1339] = in[173] | in[217]; 
    assign layer_0[1340] = in[56] | in[62]; 
    assign layer_0[1341] = ~in[134] | (in[134] & in[140]); 
    assign layer_0[1342] = in[251] | in[203]; 
    assign layer_0[1343] = in[212] & ~in[105]; 
    assign layer_0[1344] = in[5] ^ in[6]; 
    assign layer_0[1345] = ~(in[89] | in[81]); 
    assign layer_0[1346] = in[167] & ~in[217]; 
    assign layer_0[1347] = in[52] ^ in[82]; 
    assign layer_0[1348] = in[101] ^ in[180]; 
    assign layer_0[1349] = ~(in[186] | in[203]); 
    assign layer_0[1350] = in[171] ^ in[203]; 
    assign layer_0[1351] = ~(in[150] | in[35]); 
    assign layer_0[1352] = ~(in[74] ^ in[76]); 
    assign layer_0[1353] = in[99] | in[164]; 
    assign layer_0[1354] = ~in[45] | (in[92] & in[45]); 
    assign layer_0[1355] = in[244]; 
    assign layer_0[1356] = ~(in[149] ^ in[166]); 
    assign layer_0[1357] = in[198] ^ in[200]; 
    assign layer_0[1358] = in[36] | in[63]; 
    assign layer_0[1359] = in[139] ^ in[141]; 
    assign layer_0[1360] = ~(in[213] ^ in[143]); 
    assign layer_0[1361] = ~(in[231] | in[71]); 
    assign layer_0[1362] = ~in[134] | (in[134] & in[85]); 
    assign layer_0[1363] = in[78] | in[212]; 
    assign layer_0[1364] = in[23] | in[227]; 
    assign layer_0[1365] = in[165] ^ in[87]; 
    assign layer_0[1366] = ~(in[107] ^ in[89]); 
    assign layer_0[1367] = in[100] ^ in[87]; 
    assign layer_0[1368] = ~(in[97] | in[28]); 
    assign layer_0[1369] = ~(in[73] ^ in[113]); 
    assign layer_0[1370] = in[76] & ~in[29]; 
    assign layer_0[1371] = ~(in[124] | in[20]); 
    assign layer_0[1372] = in[93] ^ in[95]; 
    assign layer_0[1373] = in[156] ^ in[92]; 
    assign layer_0[1374] = in[236] ^ in[248]; 
    assign layer_0[1375] = in[164] ^ in[162]; 
    assign layer_0[1376] = in[134] | in[210]; 
    assign layer_0[1377] = ~(in[66] | in[70]); 
    assign layer_0[1378] = ~(in[120] ^ in[91]); 
    assign layer_0[1379] = ~(in[5] | in[7]); 
    assign layer_0[1380] = ~(in[230] ^ in[236]); 
    assign layer_0[1381] = in[159] ^ in[42]; 
    assign layer_0[1382] = ~in[76] | (in[122] & in[76]); 
    assign layer_0[1383] = ~(in[154] | in[46]); 
    assign layer_0[1384] = ~(in[63] | in[243]); 
    assign layer_0[1385] = in[71]; 
    assign layer_0[1386] = in[218] & ~in[109]; 
    assign layer_0[1387] = in[47] | in[95]; 
    assign layer_0[1388] = in[216] & in[214]; 
    assign layer_0[1389] = in[168] & ~in[133]; 
    assign layer_0[1390] = ~(in[136] | in[9]); 
    assign layer_0[1391] = ~in[151] | (in[151] & in[98]); 
    assign layer_0[1392] = in[154] & in[184]; 
    assign layer_0[1393] = in[26] ^ in[28]; 
    assign layer_0[1394] = in[214] | in[125]; 
    assign layer_0[1395] = ~(in[214] ^ in[182]); 
    assign layer_0[1396] = in[152] ^ in[105]; 
    assign layer_0[1397] = in[87] ^ in[67]; 
    assign layer_0[1398] = in[94] ^ in[77]; 
    assign layer_0[1399] = ~(in[153] ^ in[83]); 
    assign layer_0[1400] = in[196] ^ in[72]; 
    assign layer_0[1401] = in[37] ^ in[54]; 
    assign layer_0[1402] = in[85] | in[83]; 
    assign layer_0[1403] = ~(in[219] ^ in[173]); 
    assign layer_0[1404] = in[173] ^ in[204]; 
    assign layer_0[1405] = ~in[120] | (in[120] & in[124]); 
    assign layer_0[1406] = ~(in[109] ^ in[84]); 
    assign layer_0[1407] = in[72] ^ in[74]; 
    assign layer_0[1408] = ~(in[71] | in[39]); 
    assign layer_0[1409] = ~(in[138] | in[24]); 
    assign layer_0[1410] = ~in[135] | (in[179] & in[135]); 
    assign layer_0[1411] = in[153] ^ in[101]; 
    assign layer_0[1412] = ~in[73] | (in[45] & in[73]); 
    assign layer_0[1413] = in[198]; 
    assign layer_0[1414] = ~in[136] | (in[136] & in[157]); 
    assign layer_0[1415] = in[154] & ~in[30]; 
    assign layer_0[1416] = in[150] ^ in[131]; 
    assign layer_0[1417] = ~in[149]; 
    assign layer_0[1418] = ~in[234]; 
    assign layer_0[1419] = ~in[218] | (in[218] & in[103]); 
    assign layer_0[1420] = ~(in[235] ^ in[92]); 
    assign layer_0[1421] = in[214] ^ in[142]; 
    assign layer_0[1422] = in[117] ^ in[103]; 
    assign layer_0[1423] = in[159] | in[171]; 
    assign layer_0[1424] = in[102] | in[130]; 
    assign layer_0[1425] = ~in[165]; 
    assign layer_0[1426] = in[131] & ~in[246]; 
    assign layer_0[1427] = ~(in[91] ^ in[88]); 
    assign layer_0[1428] = ~(in[173] ^ in[171]); 
    assign layer_0[1429] = in[73]; 
    assign layer_0[1430] = in[124] | in[45]; 
    assign layer_0[1431] = ~in[102] | (in[187] & in[102]); 
    assign layer_0[1432] = ~(in[207] ^ in[104]); 
    assign layer_0[1433] = ~in[110]; 
    assign layer_0[1434] = in[139] & ~in[214]; 
    assign layer_0[1435] = in[183] ^ in[181]; 
    assign layer_0[1436] = ~(in[130] ^ in[132]); 
    assign layer_0[1437] = ~(in[41] ^ in[251]); 
    assign layer_0[1438] = ~(in[233] ^ in[117]); 
    assign layer_0[1439] = in[104]; 
    assign layer_0[1440] = in[143] | in[50]; 
    assign layer_0[1441] = in[164] | in[67]; 
    assign layer_0[1442] = in[62] | in[28]; 
    assign layer_0[1443] = in[117] ^ in[130]; 
    assign layer_0[1444] = ~(in[70] ^ in[38]); 
    assign layer_0[1445] = ~(in[40] ^ in[164]); 
    assign layer_0[1446] = in[132] ^ in[134]; 
    assign layer_0[1447] = ~(in[115] ^ in[132]); 
    assign layer_0[1448] = in[153] ^ in[122]; 
    assign layer_0[1449] = in[42] & ~in[62]; 
    assign layer_0[1450] = ~(in[137] ^ in[182]); 
    assign layer_0[1451] = ~(in[60] | in[61]); 
    assign layer_0[1452] = ~in[200] | (in[235] & in[200]); 
    assign layer_0[1453] = ~in[69]; 
    assign layer_0[1454] = in[216] & ~in[210]; 
    assign layer_0[1455] = in[69] & ~in[171]; 
    assign layer_0[1456] = in[163] ^ in[135]; 
    assign layer_0[1457] = in[78] ^ in[90]; 
    assign layer_0[1458] = ~(in[139] | in[110]); 
    assign layer_0[1459] = ~(in[49] | in[168]); 
    assign layer_0[1460] = ~(in[243] | in[146]); 
    assign layer_0[1461] = ~(in[59] | in[139]); 
    assign layer_0[1462] = in[217] ^ in[37]; 
    assign layer_0[1463] = ~(in[118] | in[237]); 
    assign layer_0[1464] = ~(in[24] | in[104]); 
    assign layer_0[1465] = in[102] ^ in[170]; 
    assign layer_0[1466] = in[60]; 
    assign layer_0[1467] = in[22]; 
    assign layer_0[1468] = in[58] | in[88]; 
    assign layer_0[1469] = in[88] & ~in[196]; 
    assign layer_0[1470] = in[54] ^ in[86]; 
    assign layer_0[1471] = in[39]; 
    assign layer_0[1472] = ~(in[88] ^ in[142]); 
    assign layer_0[1473] = in[132] ^ in[151]; 
    assign layer_0[1474] = in[5] & ~in[162]; 
    assign layer_0[1475] = ~(in[93] ^ in[55]); 
    assign layer_0[1476] = in[187]; 
    assign layer_0[1477] = ~(in[53] | in[90]); 
    assign layer_0[1478] = ~(in[247] | in[214]); 
    assign layer_0[1479] = ~in[197] | (in[197] & in[149]); 
    assign layer_0[1480] = in[154] ^ in[53]; 
    assign layer_0[1481] = ~(in[87] ^ in[55]); 
    assign layer_0[1482] = in[193] ^ in[157]; 
    assign layer_0[1483] = in[166] | in[151]; 
    assign layer_0[1484] = ~(in[131] | in[133]); 
    assign layer_0[1485] = in[228]; 
    assign layer_0[1486] = in[115] & ~in[228]; 
    assign layer_0[1487] = ~in[188] | (in[207] & in[188]); 
    assign layer_0[1488] = ~(in[68] ^ in[120]); 
    assign layer_0[1489] = ~(in[195] | in[214]); 
    assign layer_0[1490] = ~(in[98] | in[148]); 
    assign layer_0[1491] = in[211] ^ in[233]; 
    assign layer_0[1492] = ~(in[134] ^ in[126]); 
    assign layer_0[1493] = ~(in[26] | in[162]); 
    assign layer_0[1494] = ~in[87]; 
    assign layer_0[1495] = in[27] ^ in[57]; 
    assign layer_0[1496] = in[136] | in[215]; 
    assign layer_0[1497] = in[196]; 
    assign layer_0[1498] = in[147] ^ in[117]; 
    assign layer_0[1499] = ~in[154] | (in[154] & in[228]); 
    assign layer_0[1500] = in[130] | in[145]; 
    assign layer_0[1501] = ~(in[7] | in[188]); 
    assign layer_0[1502] = ~(in[132] ^ in[83]); 
    assign layer_0[1503] = ~(in[194] | in[210]); 
    assign layer_0[1504] = in[39] ^ in[87]; 
    assign layer_0[1505] = ~(in[41] ^ in[99]); 
    assign layer_0[1506] = in[119] ^ in[133]; 
    assign layer_0[1507] = ~(in[244] ^ in[155]); 
    assign layer_0[1508] = in[92] ^ in[199]; 
    assign layer_0[1509] = ~(in[162] ^ in[122]); 
    assign layer_0[1510] = in[133] | in[251]; 
    assign layer_0[1511] = ~(in[60] ^ in[103]); 
    assign layer_0[1512] = ~(in[152] | in[108]); 
    assign layer_0[1513] = in[22] & ~in[242]; 
    assign layer_0[1514] = ~(in[43] ^ in[75]); 
    assign layer_0[1515] = ~(in[56] & in[85]); 
    assign layer_0[1516] = in[99] ^ in[85]; 
    assign layer_0[1517] = in[95]; 
    assign layer_0[1518] = in[59] & ~in[9]; 
    assign layer_0[1519] = ~(in[164] ^ in[133]); 
    assign layer_0[1520] = in[178] ^ in[180]; 
    assign layer_0[1521] = in[146] & ~in[236]; 
    assign layer_0[1522] = in[156] ^ in[142]; 
    assign layer_0[1523] = ~(in[126] | in[125]); 
    assign layer_0[1524] = in[79] & ~in[100]; 
    assign layer_0[1525] = in[107] ^ in[124]; 
    assign layer_0[1526] = ~in[205]; 
    assign layer_0[1527] = ~in[146]; 
    assign layer_0[1528] = in[150] & ~in[78]; 
    assign layer_0[1529] = in[146] | in[67]; 
    assign layer_0[1530] = ~(in[98] | in[78]); 
    assign layer_0[1531] = ~in[156]; 
    assign layer_0[1532] = ~in[166]; 
    assign layer_0[1533] = in[76] & ~in[217]; 
    assign layer_0[1534] = ~(in[230] | in[246]); 
    assign layer_0[1535] = in[41] ^ in[84]; 
    assign layer_0[1536] = in[120] | in[231]; 
    assign layer_0[1537] = ~(in[245] ^ in[197]); 
    assign layer_0[1538] = in[119] & ~in[70]; 
    assign layer_0[1539] = in[100] & ~in[155]; 
    assign layer_0[1540] = ~(in[230] ^ in[215]); 
    assign layer_0[1541] = ~in[151] | (in[151] & in[217]); 
    assign layer_0[1542] = ~(in[84] | in[135]); 
    assign layer_0[1543] = in[202] | in[202]; 
    assign layer_0[1544] = ~in[107] | (in[220] & in[107]); 
    assign layer_0[1545] = ~(in[134] ^ in[126]); 
    assign layer_0[1546] = ~in[150]; 
    assign layer_0[1547] = ~(in[87] | in[120]); 
    assign layer_0[1548] = ~(in[196] | in[183]); 
    assign layer_0[1549] = in[137]; 
    assign layer_0[1550] = ~(in[6] | in[84]); 
    assign layer_0[1551] = ~(in[189] ^ in[157]); 
    assign layer_0[1552] = in[8]; 
    assign layer_0[1553] = ~(in[211] | in[222]); 
    assign layer_0[1554] = in[221] & ~in[125]; 
    assign layer_0[1555] = in[95] ^ in[174]; 
    assign layer_0[1556] = in[25] ^ in[57]; 
    assign layer_0[1557] = in[215] | in[197]; 
    assign layer_0[1558] = ~(in[21] | in[50]); 
    assign layer_0[1559] = in[8] ^ in[10]; 
    assign layer_0[1560] = in[41] ^ in[73]; 
    assign layer_0[1561] = ~(in[151] & in[148]); 
    assign layer_0[1562] = ~(in[149] ^ in[127]); 
    assign layer_0[1563] = in[43] | in[58]; 
    assign layer_0[1564] = in[182] & ~in[249]; 
    assign layer_0[1565] = ~(in[77] ^ in[198]); 
    assign layer_0[1566] = ~(in[65] | in[34]); 
    assign layer_0[1567] = in[230] & ~in[183]; 
    assign layer_0[1568] = ~(in[83] | in[212]); 
    assign layer_0[1569] = in[84] ^ in[133]; 
    assign layer_0[1570] = ~in[40] | (in[40] & in[140]); 
    assign layer_0[1571] = ~(in[103] ^ in[134]); 
    assign layer_0[1572] = ~in[163] | (in[250] & in[163]); 
    assign layer_0[1573] = in[248]; 
    assign layer_0[1574] = ~(in[164] | in[84]); 
    assign layer_0[1575] = in[120] & ~in[171]; 
    assign layer_0[1576] = ~(in[183] ^ in[98]); 
    assign layer_0[1577] = ~(in[165] ^ in[202]); 
    assign layer_0[1578] = ~(in[150] | in[134]); 
    assign layer_0[1579] = in[181]; 
    assign layer_0[1580] = ~(in[116] ^ in[102]); 
    assign layer_0[1581] = in[136]; 
    assign layer_0[1582] = in[127] | in[110]; 
    assign layer_0[1583] = in[73] ^ in[75]; 
    assign layer_0[1584] = ~(in[45] ^ in[226]); 
    assign layer_0[1585] = in[168] ^ in[121]; 
    assign layer_0[1586] = in[11] & ~in[78]; 
    assign layer_0[1587] = in[68] ^ in[70]; 
    assign layer_0[1588] = ~(in[83] | in[85]); 
    assign layer_0[1589] = in[168] | in[137]; 
    assign layer_0[1590] = in[51] | in[178]; 
    assign layer_0[1591] = in[119] & ~in[52]; 
    assign layer_0[1592] = ~in[72]; 
    assign layer_0[1593] = ~(in[27] ^ in[56]); 
    assign layer_0[1594] = in[90] | in[203]; 
    assign layer_0[1595] = ~(in[79] ^ in[183]); 
    assign layer_0[1596] = ~(in[24] ^ in[71]); 
    assign layer_0[1597] = ~(in[78] ^ in[51]); 
    assign layer_0[1598] = in[135] ^ in[120]; 
    assign layer_0[1599] = ~(in[56] ^ in[95]); 
    assign layer_0[1600] = in[167] & ~in[63]; 
    assign layer_0[1601] = in[163]; 
    assign layer_0[1602] = ~(in[167] & in[137]); 
    assign layer_0[1603] = ~(in[61] ^ in[75]); 
    assign layer_0[1604] = in[46]; 
    assign layer_0[1605] = in[78] | in[76]; 
    assign layer_0[1606] = in[17] & in[253]; 
    assign layer_0[1607] = in[164] ^ in[146]; 
    assign layer_0[1608] = in[37] ^ in[52]; 
    assign layer_0[1609] = in[229] ^ in[198]; 
    assign layer_0[1610] = in[150] | in[114]; 
    assign layer_0[1611] = ~(in[140] ^ in[171]); 
    assign layer_0[1612] = in[47] | in[79]; 
    assign layer_0[1613] = ~(in[146] | in[109]); 
    assign layer_0[1614] = in[104]; 
    assign layer_0[1615] = ~(in[117] ^ in[115]); 
    assign layer_0[1616] = ~(in[140] ^ in[136]); 
    assign layer_0[1617] = in[198] ^ in[248]; 
    assign layer_0[1618] = ~in[82] | (in[197] & in[82]); 
    assign layer_0[1619] = in[164] ^ in[183]; 
    assign layer_0[1620] = in[155] & ~in[35]; 
    assign layer_0[1621] = in[146] ^ in[133]; 
    assign layer_0[1622] = ~(in[102] ^ in[78]); 
    assign layer_0[1623] = in[90] | in[107]; 
    assign layer_0[1624] = ~in[185]; 
    assign layer_0[1625] = ~(in[100] ^ in[102]); 
    assign layer_0[1626] = in[83] ^ in[245]; 
    assign layer_0[1627] = ~in[120] | (in[109] & in[120]); 
    assign layer_0[1628] = in[140] ^ in[123]; 
    assign layer_0[1629] = in[165] ^ in[163]; 
    assign layer_0[1630] = in[119] & ~in[101]; 
    assign layer_0[1631] = in[216] & ~in[169]; 
    assign layer_0[1632] = ~in[148]; 
    assign layer_0[1633] = in[146] ^ in[196]; 
    assign layer_0[1634] = in[153] & ~in[74]; 
    assign layer_0[1635] = ~(in[164] ^ in[150]); 
    assign layer_0[1636] = in[133] ^ in[115]; 
    assign layer_0[1637] = ~in[59] | (in[220] & in[59]); 
    assign layer_0[1638] = ~(in[44] ^ in[76]); 
    assign layer_0[1639] = ~in[153] | (in[153] & in[21]); 
    assign layer_0[1640] = in[23] ^ in[58]; 
    assign layer_0[1641] = in[251] | in[137]; 
    assign layer_0[1642] = in[210]; 
    assign layer_0[1643] = ~(in[102] ^ in[35]); 
    assign layer_0[1644] = ~in[214]; 
    assign layer_0[1645] = ~in[78]; 
    assign layer_0[1646] = ~(in[27] | in[184]); 
    assign layer_0[1647] = ~(in[231] ^ in[243]); 
    assign layer_0[1648] = ~in[42]; 
    assign layer_0[1649] = ~in[133] | (in[133] & in[188]); 
    assign layer_0[1650] = ~in[77]; 
    assign layer_0[1651] = in[120]; 
    assign layer_0[1652] = ~(in[163] | in[117]); 
    assign layer_0[1653] = ~in[59]; 
    assign layer_0[1654] = in[152] | in[23]; 
    assign layer_0[1655] = in[113] | in[110]; 
    assign layer_0[1656] = ~(in[83] ^ in[35]); 
    assign layer_0[1657] = ~(in[140] | in[173]); 
    assign layer_0[1658] = in[81] | in[66]; 
    assign layer_0[1659] = in[104]; 
    assign layer_0[1660] = ~in[122] | (in[109] & in[122]); 
    assign layer_0[1661] = in[72] | in[71]; 
    assign layer_0[1662] = in[57] ^ in[156]; 
    assign layer_0[1663] = in[72]; 
    assign layer_0[1664] = in[183] | in[183]; 
    assign layer_0[1665] = in[230] & ~in[187]; 
    assign layer_0[1666] = in[134] & ~in[113]; 
    assign layer_0[1667] = in[44] | in[27]; 
    assign layer_0[1668] = ~(in[196] ^ in[204]); 
    assign layer_0[1669] = in[23] ^ in[26]; 
    assign layer_0[1670] = in[69] ^ in[37]; 
    assign layer_0[1671] = ~(in[146] | in[134]); 
    assign layer_0[1672] = in[121] ^ in[178]; 
    assign layer_0[1673] = in[166] | in[104]; 
    assign layer_0[1674] = in[54] ^ in[60]; 
    assign layer_0[1675] = in[69] ^ in[23]; 
    assign layer_0[1676] = ~(in[55] ^ in[23]); 
    assign layer_0[1677] = ~(in[119] | in[77]); 
    assign layer_0[1678] = in[212] | in[210]; 
    assign layer_0[1679] = ~in[44] | (in[195] & in[44]); 
    assign layer_0[1680] = ~(in[72] ^ in[126]); 
    assign layer_0[1681] = in[57] | in[41]; 
    assign layer_0[1682] = in[55] ^ in[9]; 
    assign layer_0[1683] = ~(in[218] ^ in[211]); 
    assign layer_0[1684] = in[58] ^ in[89]; 
    assign layer_0[1685] = in[125]; 
    assign layer_0[1686] = in[180] | in[135]; 
    assign layer_0[1687] = ~(in[53] ^ in[92]); 
    assign layer_0[1688] = in[93]; 
    assign layer_0[1689] = in[136] | in[104]; 
    assign layer_0[1690] = ~(in[130] ^ in[116]); 
    assign layer_0[1691] = ~in[106] | (in[106] & in[5]); 
    assign layer_0[1692] = in[146] ^ in[62]; 
    assign layer_0[1693] = in[74] & ~in[71]; 
    assign layer_0[1694] = in[130] ^ in[129]; 
    assign layer_0[1695] = in[74] ^ in[125]; 
    assign layer_0[1696] = ~in[198] | (in[27] & in[198]); 
    assign layer_0[1697] = ~(in[62] | in[163]); 
    assign layer_0[1698] = in[102] | in[93]; 
    assign layer_0[1699] = in[158] | in[139]; 
    assign layer_0[1700] = ~(in[231] | in[179]); 
    assign layer_0[1701] = in[81] | in[66]; 
    assign layer_0[1702] = in[233]; 
    assign layer_0[1703] = in[181]; 
    assign layer_0[1704] = in[182] & ~in[115]; 
    assign layer_0[1705] = ~(in[248] ^ in[21]); 
    assign layer_0[1706] = in[120] ^ in[104]; 
    assign layer_0[1707] = in[103] | in[132]; 
    assign layer_0[1708] = ~(in[21] ^ in[8]); 
    assign layer_0[1709] = ~(in[37] | in[26]); 
    assign layer_0[1710] = in[126]; 
    assign layer_0[1711] = in[63] ^ in[241]; 
    assign layer_0[1712] = ~(in[102] | in[117]); 
    assign layer_0[1713] = in[70] & ~in[183]; 
    assign layer_0[1714] = in[56]; 
    assign layer_0[1715] = ~in[199] | (in[58] & in[199]); 
    assign layer_0[1716] = in[149] & ~in[73]; 
    assign layer_0[1717] = ~in[200] | (in[69] & in[200]); 
    assign layer_0[1718] = ~in[140] | (in[180] & in[140]); 
    assign layer_0[1719] = in[59] & ~in[25]; 
    assign layer_0[1720] = in[84] ^ in[118]; 
    assign layer_0[1721] = in[135] ^ in[103]; 
    assign layer_0[1722] = in[120] | in[151]; 
    assign layer_0[1723] = in[22] ^ in[136]; 
    assign layer_0[1724] = ~(in[60] | in[143]); 
    assign layer_0[1725] = in[177]; 
    assign layer_0[1726] = in[165] ^ in[167]; 
    assign layer_0[1727] = ~(in[119] ^ in[148]); 
    assign layer_0[1728] = ~in[105] | (in[156] & in[105]); 
    assign layer_0[1729] = in[137] | in[13]; 
    assign layer_0[1730] = ~in[59] | (in[59] & in[44]); 
    assign layer_0[1731] = ~(in[153] ^ in[114]); 
    assign layer_0[1732] = in[78] ^ in[56]; 
    assign layer_0[1733] = ~(in[74] | in[156]); 
    assign layer_0[1734] = ~in[87] | (in[179] & in[87]); 
    assign layer_0[1735] = ~(in[173] ^ in[195]); 
    assign layer_0[1736] = in[164] ^ in[181]; 
    assign layer_0[1737] = ~in[104]; 
    assign layer_0[1738] = ~(in[161] | in[200]); 
    assign layer_0[1739] = ~(in[34] | in[6]); 
    assign layer_0[1740] = ~(in[86] ^ in[170]); 
    assign layer_0[1741] = in[195] ^ in[220]; 
    assign layer_0[1742] = ~(in[214] ^ in[245]); 
    assign layer_0[1743] = ~in[170] | (in[142] & in[170]); 
    assign layer_0[1744] = in[38] | in[21]; 
    assign layer_0[1745] = ~(in[166] | in[250]); 
    assign layer_0[1746] = ~in[245] | (in[245] & in[212]); 
    assign layer_0[1747] = ~(in[52] ^ in[85]); 
    assign layer_0[1748] = ~in[44] | (in[122] & in[44]); 
    assign layer_0[1749] = in[154] ^ in[21]; 
    assign layer_0[1750] = ~(in[100] ^ in[132]); 
    assign layer_0[1751] = in[70] ^ in[39]; 
    assign layer_0[1752] = ~in[183]; 
    assign layer_0[1753] = ~(in[119] ^ in[113]); 
    assign layer_0[1754] = ~(in[77] | in[89]); 
    assign layer_0[1755] = in[61] ^ in[95]; 
    assign layer_0[1756] = ~(in[47] | in[53]); 
    assign layer_0[1757] = in[212] & ~in[123]; 
    assign layer_0[1758] = in[104] & ~in[118]; 
    assign layer_0[1759] = in[7] ^ in[213]; 
    assign layer_0[1760] = ~(in[173] ^ in[41]); 
    assign layer_0[1761] = in[138]; 
    assign layer_0[1762] = ~(in[148] ^ in[130]); 
    assign layer_0[1763] = in[170] | in[155]; 
    assign layer_0[1764] = in[70] ^ in[24]; 
    assign layer_0[1765] = ~(in[172] | in[197]); 
    assign layer_0[1766] = ~(in[153] | in[135]); 
    assign layer_0[1767] = ~(in[116] ^ in[113]); 
    assign layer_0[1768] = in[12] | in[30]; 
    assign layer_0[1769] = in[131] | in[20]; 
    assign layer_0[1770] = in[210] | in[88]; 
    assign layer_0[1771] = in[137]; 
    assign layer_0[1772] = ~in[104]; 
    assign layer_0[1773] = ~(in[165] ^ in[167]); 
    assign layer_0[1774] = in[78] ^ in[91]; 
    assign layer_0[1775] = ~(in[249] ^ in[220]); 
    assign layer_0[1776] = in[249] ^ in[235]; 
    assign layer_0[1777] = ~(in[198] | in[196]); 
    assign layer_0[1778] = in[20] ^ in[170]; 
    assign layer_0[1779] = in[169] ^ in[195]; 
    assign layer_0[1780] = in[218] | in[167]; 
    assign layer_0[1781] = in[181] ^ in[150]; 
    assign layer_0[1782] = ~(in[59] | in[74]); 
    assign layer_0[1783] = in[123]; 
    assign layer_0[1784] = ~(in[99] ^ in[121]); 
    assign layer_0[1785] = in[125] | in[86]; 
    assign layer_0[1786] = ~(in[85] | in[83]); 
    assign layer_0[1787] = in[157]; 
    assign layer_0[1788] = ~(in[42] ^ in[89]); 
    assign layer_0[1789] = in[221] ^ in[106]; 
    assign layer_0[1790] = in[83]; 
    assign layer_0[1791] = ~(in[76] ^ in[123]); 
    assign layer_0[1792] = ~in[244] | (in[41] & in[244]); 
    assign layer_0[1793] = ~(in[91] ^ in[94]); 
    assign layer_0[1794] = in[248] ^ in[219]; 
    assign layer_0[1795] = ~(in[253] ^ in[235]); 
    assign layer_0[1796] = ~(in[183] ^ in[100]); 
    assign layer_0[1797] = ~(in[46] ^ in[29]); 
    assign layer_0[1798] = ~(in[151] ^ in[27]); 
    assign layer_0[1799] = in[163] ^ in[180]; 
    assign layer_0[1800] = ~(in[116] | in[92]); 
    assign layer_0[1801] = in[68] ^ in[82]; 
    assign layer_0[1802] = in[75] & ~in[87]; 
    assign layer_0[1803] = in[157] | in[75]; 
    assign layer_0[1804] = ~in[41] | (in[180] & in[41]); 
    assign layer_0[1805] = ~(in[84] ^ in[67]); 
    assign layer_0[1806] = ~(in[52] ^ in[41]); 
    assign layer_0[1807] = in[136] & ~in[95]; 
    assign layer_0[1808] = in[71] ^ in[175]; 
    assign layer_0[1809] = in[142] ^ in[157]; 
    assign layer_0[1810] = ~(in[88] ^ in[214]); 
    assign layer_0[1811] = in[177] | in[243]; 
    assign layer_0[1812] = in[53] ^ in[86]; 
    assign layer_0[1813] = in[54] ^ in[7]; 
    assign layer_0[1814] = in[56] | in[86]; 
    assign layer_0[1815] = in[170] | in[27]; 
    assign layer_0[1816] = ~(in[63] ^ in[30]); 
    assign layer_0[1817] = in[215]; 
    assign layer_0[1818] = in[26] ^ in[75]; 
    assign layer_0[1819] = in[84] ^ in[70]; 
    assign layer_0[1820] = in[198] & in[168]; 
    assign layer_0[1821] = in[120] & ~in[53]; 
    assign layer_0[1822] = ~(in[27] ^ in[194]); 
    assign layer_0[1823] = ~(in[50] ^ in[92]); 
    assign layer_0[1824] = ~(in[123] | in[98]); 
    assign layer_0[1825] = in[150] & ~in[157]; 
    assign layer_0[1826] = in[195] | in[40]; 
    assign layer_0[1827] = in[174] ^ in[206]; 
    assign layer_0[1828] = in[106] ^ in[248]; 
    assign layer_0[1829] = ~in[213]; 
    assign layer_0[1830] = in[121]; 
    assign layer_0[1831] = ~in[73] | (in[235] & in[73]); 
    assign layer_0[1832] = in[71] ^ in[37]; 
    assign layer_0[1833] = ~(in[200] ^ in[232]); 
    assign layer_0[1834] = ~in[181] | (in[244] & in[181]); 
    assign layer_0[1835] = in[135] & ~in[155]; 
    assign layer_0[1836] = ~(in[76] ^ in[106]); 
    assign layer_0[1837] = in[199] ^ in[44]; 
    assign layer_0[1838] = ~in[125] | (in[125] & in[73]); 
    assign layer_0[1839] = ~(in[38] ^ in[232]); 
    assign layer_0[1840] = in[162] & ~in[210]; 
    assign layer_0[1841] = in[251] & ~in[171]; 
    assign layer_0[1842] = in[181] | in[221]; 
    assign layer_0[1843] = in[81] | in[52]; 
    assign layer_0[1844] = in[53]; 
    assign layer_0[1845] = in[105] ^ in[167]; 
    assign layer_0[1846] = in[92] ^ in[123]; 
    assign layer_0[1847] = in[216] ^ in[248]; 
    assign layer_0[1848] = in[236] ^ in[205]; 
    assign layer_0[1849] = ~(in[167] | in[121]); 
    assign layer_0[1850] = in[214] ^ in[167]; 
    assign layer_0[1851] = in[199] | in[198]; 
    assign layer_0[1852] = in[135] & ~in[164]; 
    assign layer_0[1853] = ~(in[60] ^ in[184]); 
    assign layer_0[1854] = ~(in[233] ^ in[246]); 
    assign layer_0[1855] = in[105] ^ in[152]; 
    assign layer_0[1856] = in[212] ^ in[71]; 
    assign layer_0[1857] = ~(in[34] ^ in[210]); 
    assign layer_0[1858] = ~in[170] | (in[221] & in[170]); 
    assign layer_0[1859] = in[212] & ~in[100]; 
    assign layer_0[1860] = ~(in[28] ^ in[194]); 
    assign layer_0[1861] = ~(in[102] ^ in[55]); 
    assign layer_0[1862] = in[182] | in[183]; 
    assign layer_0[1863] = ~in[182] | (in[182] & in[61]); 
    assign layer_0[1864] = ~in[231]; 
    assign layer_0[1865] = in[216] & ~in[147]; 
    assign layer_0[1866] = ~(in[91] ^ in[62]); 
    assign layer_0[1867] = ~in[154] | (in[154] & in[126]); 
    assign layer_0[1868] = ~(in[155] ^ in[170]); 
    assign layer_0[1869] = ~(in[24] ^ in[44]); 
    assign layer_0[1870] = ~(in[212] | in[201]); 
    assign layer_0[1871] = ~(in[236] | in[41]); 
    assign layer_0[1872] = ~(in[180] | in[202]); 
    assign layer_0[1873] = ~(in[219] ^ in[172]); 
    assign layer_0[1874] = in[24] ^ in[56]; 
    assign layer_0[1875] = in[37] | in[90]; 
    assign layer_0[1876] = in[43]; 
    assign layer_0[1877] = in[168] ^ in[150]; 
    assign layer_0[1878] = in[75] | in[76]; 
    assign layer_0[1879] = in[104] & ~in[186]; 
    assign layer_0[1880] = in[212] ^ in[166]; 
    assign layer_0[1881] = ~in[140] | (in[212] & in[140]); 
    assign layer_0[1882] = ~(in[163] ^ in[132]); 
    assign layer_0[1883] = ~(in[168] | in[94]); 
    assign layer_0[1884] = ~(in[77] ^ in[109]); 
    assign layer_0[1885] = in[186] & ~in[131]; 
    assign layer_0[1886] = in[138] ^ in[106]; 
    assign layer_0[1887] = ~in[122] | (in[122] & in[228]); 
    assign layer_0[1888] = in[201] | in[21]; 
    assign layer_0[1889] = ~(in[44] ^ in[75]); 
    assign layer_0[1890] = in[248] ^ in[202]; 
    assign layer_0[1891] = in[72] & ~in[60]; 
    assign layer_0[1892] = in[200] & ~in[79]; 
    assign layer_0[1893] = ~(in[166] ^ in[247]); 
    assign layer_0[1894] = in[236] ^ in[249]; 
    assign layer_0[1895] = ~in[245]; 
    assign layer_0[1896] = ~(in[211] ^ in[226]); 
    assign layer_0[1897] = in[200] ^ in[166]; 
    assign layer_0[1898] = ~(in[191] ^ in[143]); 
    assign layer_0[1899] = in[102] & ~in[59]; 
    assign layer_0[1900] = ~(in[219] ^ in[182]); 
    assign layer_0[1901] = ~(in[184] | in[206]); 
    assign layer_0[1902] = ~(in[167] | in[135]); 
    assign layer_0[1903] = ~(in[125] | in[127]); 
    assign layer_0[1904] = ~(in[102] ^ in[251]); 
    assign layer_0[1905] = in[147] | in[76]; 
    assign layer_0[1906] = in[194] ^ in[213]; 
    assign layer_0[1907] = ~(in[93] | in[36]); 
    assign layer_0[1908] = ~in[170] | (in[120] & in[170]); 
    assign layer_0[1909] = ~in[57] | (in[57] & in[121]); 
    assign layer_0[1910] = ~(in[153] ^ in[120]); 
    assign layer_0[1911] = ~(in[21] | in[237]); 
    assign layer_0[1912] = ~(in[9] ^ in[12]); 
    assign layer_0[1913] = ~in[232] | (in[232] & in[19]); 
    assign layer_0[1914] = in[118] ^ in[104]; 
    assign layer_0[1915] = in[12] & ~in[54]; 
    assign layer_0[1916] = in[172] & ~in[254]; 
    assign layer_0[1917] = ~(in[71] ^ in[157]); 
    assign layer_0[1918] = ~(in[81] | in[200]); 
    assign layer_0[1919] = in[149] | in[148]; 
    assign layer_0[1920] = in[242] ^ in[86]; 
    assign layer_0[1921] = ~(in[215] ^ in[246]); 
    assign layer_0[1922] = in[184] ^ in[46]; 
    assign layer_0[1923] = ~(in[98] ^ in[100]); 
    assign layer_0[1924] = in[114] ^ in[101]; 
    assign layer_0[1925] = ~(in[203] ^ in[201]); 
    assign layer_0[1926] = in[7]; 
    assign layer_0[1927] = ~(in[244] ^ in[62]); 
    assign layer_0[1928] = ~in[66]; 
    assign layer_0[1929] = in[117] | in[115]; 
    assign layer_0[1930] = ~(in[34] ^ in[60]); 
    assign layer_0[1931] = in[105] | in[92]; 
    assign layer_0[1932] = in[75]; 
    assign layer_0[1933] = in[121] & ~in[203]; 
    assign layer_0[1934] = in[149] | in[133]; 
    assign layer_0[1935] = ~(in[229] | in[53]); 
    assign layer_0[1936] = in[75] ^ in[44]; 
    assign layer_0[1937] = ~(in[250] | in[163]); 
    assign layer_0[1938] = ~in[163] | (in[163] & in[122]); 
    assign layer_0[1939] = in[58] & ~in[38]; 
    assign layer_0[1940] = in[97] ^ in[119]; 
    assign layer_0[1941] = ~(in[100] ^ in[102]); 
    assign layer_0[1942] = in[116] | in[241]; 
    assign layer_0[1943] = ~in[166]; 
    assign layer_0[1944] = ~(in[96] | in[249]); 
    assign layer_0[1945] = ~(in[235] | in[178]); 
    assign layer_0[1946] = ~(in[59] | in[141]); 
    assign layer_0[1947] = ~(in[178] ^ in[150]); 
    assign layer_0[1948] = ~in[34]; 
    assign layer_0[1949] = ~(in[54] | in[37]); 
    assign layer_0[1950] = in[165] ^ in[134]; 
    assign layer_0[1951] = ~(in[124] ^ in[250]); 
    assign layer_0[1952] = ~in[91] | (in[91] & in[104]); 
    assign layer_0[1953] = in[87] | in[181]; 
    assign layer_0[1954] = in[179] ^ in[199]; 
    assign layer_0[1955] = in[125] | in[140]; 
    assign layer_0[1956] = ~(in[172] ^ in[50]); 
    assign layer_0[1957] = in[82] ^ in[25]; 
    assign layer_0[1958] = ~(in[91] ^ in[55]); 
    assign layer_0[1959] = in[53] ^ in[85]; 
    assign layer_0[1960] = ~in[198] | (in[198] & in[141]); 
    assign layer_0[1961] = in[33] | in[12]; 
    assign layer_0[1962] = in[9] | in[85]; 
    assign layer_0[1963] = in[105] & ~in[92]; 
    assign layer_0[1964] = in[113] ^ in[41]; 
    assign layer_0[1965] = in[37] | in[107]; 
    assign layer_0[1966] = ~in[41]; 
    assign layer_0[1967] = in[35]; 
    assign layer_0[1968] = in[53] ^ in[89]; 
    assign layer_0[1969] = ~in[142] | (in[235] & in[142]); 
    assign layer_0[1970] = ~(in[180] ^ in[182]); 
    assign layer_0[1971] = in[155] ^ in[51]; 
    assign layer_0[1972] = ~(in[43] ^ in[198]); 
    assign layer_0[1973] = ~(in[221] ^ in[95]); 
    assign layer_0[1974] = in[103]; 
    assign layer_0[1975] = ~(in[186] ^ in[37]); 
    assign layer_0[1976] = ~(in[134] | in[68]); 
    assign layer_0[1977] = ~in[169] | (in[5] & in[169]); 
    assign layer_0[1978] = in[234] & ~in[166]; 
    assign layer_0[1979] = ~in[102] | (in[102] & in[73]); 
    assign layer_0[1980] = in[58] & ~in[156]; 
    assign layer_0[1981] = ~(in[140] | in[204]); 
    assign layer_0[1982] = in[40] ^ in[87]; 
    assign layer_0[1983] = ~(in[171] ^ in[152]); 
    assign layer_0[1984] = in[195] ^ in[216]; 
    assign layer_0[1985] = in[221] | in[175]; 
    assign layer_0[1986] = ~(in[243] | in[223]); 
    assign layer_0[1987] = ~(in[109] | in[84]); 
    assign layer_0[1988] = ~(in[245] | in[210]); 
    assign layer_0[1989] = in[213] & in[57]; 
    assign layer_0[1990] = ~in[90] | (in[90] & in[183]); 
    assign layer_0[1991] = in[235] ^ in[118]; 
    assign layer_0[1992] = ~in[93]; 
    assign layer_0[1993] = in[19] ^ in[92]; 
    assign layer_0[1994] = in[186] | in[140]; 
    assign layer_0[1995] = in[108] ^ in[59]; 
    assign layer_0[1996] = in[125]; 
    assign layer_0[1997] = ~in[135] | (in[135] & in[242]); 
    assign layer_0[1998] = in[52] ^ in[83]; 
    assign layer_0[1999] = ~in[199]; 
    assign layer_0[2000] = in[203] | in[30]; 
    assign layer_0[2001] = ~(in[182] | in[165]); 
    assign layer_0[2002] = in[109]; 
    assign layer_0[2003] = ~(in[51] ^ in[36]); 
    assign layer_0[2004] = ~(in[88] ^ in[118]); 
    assign layer_0[2005] = in[139] ^ in[187]; 
    assign layer_0[2006] = ~(in[9] | in[146]); 
    assign layer_0[2007] = in[86] ^ in[41]; 
    assign layer_0[2008] = in[105] & in[104]; 
    assign layer_0[2009] = in[100] ^ in[87]; 
    assign layer_0[2010] = in[36] | in[44]; 
    assign layer_0[2011] = in[68]; 
    assign layer_0[2012] = ~(in[12] ^ in[198]); 
    assign layer_0[2013] = ~(in[94] | in[174]); 
    assign layer_0[2014] = ~in[202] | (in[202] & in[146]); 
    assign layer_0[2015] = ~in[140] | (in[189] & in[140]); 
    assign layer_0[2016] = ~(in[28] ^ in[26]); 
    assign layer_0[2017] = ~(in[115] | in[163]); 
    assign layer_0[2018] = in[181] ^ in[211]; 
    assign layer_0[2019] = ~(in[227] ^ in[24]); 
    assign layer_0[2020] = ~(in[56] | in[230]); 
    assign layer_0[2021] = in[198] & ~in[107]; 
    assign layer_0[2022] = ~(in[85] ^ in[99]); 
    assign layer_0[2023] = in[124] ^ in[167]; 
    assign layer_0[2024] = in[99] ^ in[98]; 
    assign layer_0[2025] = in[51] ^ in[229]; 
    assign layer_0[2026] = ~(in[109] ^ in[140]); 
    assign layer_0[2027] = in[37] | in[150]; 
    assign layer_0[2028] = ~(in[168] ^ in[250]); 
    assign layer_0[2029] = ~in[202] | (in[198] & in[202]); 
    assign layer_0[2030] = ~in[137] | (in[137] & in[179]); 
    assign layer_0[2031] = ~(in[91] ^ in[93]); 
    assign layer_0[2032] = ~in[155] | (in[137] & in[155]); 
    assign layer_0[2033] = in[90] ^ in[59]; 
    assign layer_0[2034] = ~(in[157] | in[105]); 
    assign layer_0[2035] = ~(in[93] ^ in[125]); 
    assign layer_0[2036] = ~(in[40] ^ in[147]); 
    assign layer_0[2037] = ~(in[156] ^ in[187]); 
    assign layer_0[2038] = in[187] ^ in[235]; 
    assign layer_0[2039] = ~(in[87] ^ in[73]); 
    assign layer_0[2040] = ~(in[231] | in[215]); 
    assign layer_0[2041] = in[90] & ~in[63]; 
    assign layer_0[2042] = ~(in[70] ^ in[84]); 
    assign layer_0[2043] = in[167] & in[136]; 
    assign layer_0[2044] = in[84] ^ in[186]; 
    assign layer_0[2045] = ~(in[220] | in[181]); 
    assign layer_0[2046] = ~in[211] | (in[211] & in[88]); 
    assign layer_0[2047] = in[149] & ~in[129]; 
    assign layer_0[2048] = ~(in[103] | in[88]); 
    assign layer_0[2049] = ~(in[167] ^ in[215]); 
    assign layer_0[2050] = ~in[73] | (in[73] & in[117]); 
    assign layer_0[2051] = ~(in[212] ^ in[214]); 
    assign layer_0[2052] = ~in[117] | (in[117] & in[140]); 
    assign layer_0[2053] = in[105] ^ in[152]; 
    assign layer_0[2054] = ~(in[211] ^ in[92]); 
    assign layer_0[2055] = ~(in[86] | in[91]); 
    assign layer_0[2056] = ~(in[116] ^ in[118]); 
    assign layer_0[2057] = ~in[202] | (in[202] & in[118]); 
    assign layer_0[2058] = in[105] & ~in[23]; 
    assign layer_0[2059] = in[59] | in[74]; 
    assign layer_0[2060] = ~in[58] | (in[58] & in[167]); 
    assign layer_0[2061] = in[25] & ~in[149]; 
    assign layer_0[2062] = ~in[105]; 
    assign layer_0[2063] = ~in[185] | (in[185] & in[25]); 
    assign layer_0[2064] = in[169] ^ in[103]; 
    assign layer_0[2065] = ~(in[203] ^ in[236]); 
    assign layer_0[2066] = ~in[82]; 
    assign layer_0[2067] = in[154] ^ in[230]; 
    assign layer_0[2068] = in[46] | in[29]; 
    assign layer_0[2069] = in[99] | in[163]; 
    assign layer_0[2070] = in[142] ^ in[29]; 
    assign layer_0[2071] = in[134] ^ in[142]; 
    assign layer_0[2072] = in[42] ^ in[166]; 
    assign layer_0[2073] = ~(in[139] & in[170]); 
    assign layer_0[2074] = ~(in[164] ^ in[182]); 
    assign layer_0[2075] = ~in[116] | (in[116] & in[165]); 
    assign layer_0[2076] = in[85] ^ in[82]; 
    assign layer_0[2077] = ~(in[100] ^ in[113]); 
    assign layer_0[2078] = in[182] ^ in[180]; 
    assign layer_0[2079] = ~(in[56] ^ in[24]); 
    assign layer_0[2080] = ~in[167] | (in[132] & in[167]); 
    assign layer_0[2081] = ~(in[11] ^ in[118]); 
    assign layer_0[2082] = in[40] | in[25]; 
    assign layer_0[2083] = ~(in[148] ^ in[131]); 
    assign layer_0[2084] = in[63] | in[114]; 
    assign layer_0[2085] = ~(in[124] ^ in[103]); 
    assign layer_0[2086] = in[94] ^ in[92]; 
    assign layer_0[2087] = in[88] & in[91]; 
    assign layer_0[2088] = ~(in[139] & in[150]); 
    assign layer_0[2089] = ~(in[162] ^ in[154]); 
    assign layer_0[2090] = in[74]; 
    assign layer_0[2091] = ~(in[75] ^ in[92]); 
    assign layer_0[2092] = ~in[153] | (in[196] & in[153]); 
    assign layer_0[2093] = in[159] | in[145]; 
    assign layer_0[2094] = ~in[73] | (in[73] & in[219]); 
    assign layer_0[2095] = in[245] | in[24]; 
    assign layer_0[2096] = in[135]; 
    assign layer_0[2097] = in[137] ^ in[178]; 
    assign layer_0[2098] = ~(in[34] | in[51]); 
    assign layer_0[2099] = in[130] | in[193]; 
    assign layer_0[2100] = in[150] ^ in[142]; 
    assign layer_0[2101] = ~(in[228] | in[245]); 
    assign layer_0[2102] = ~in[183] | (in[183] & in[212]); 
    assign layer_0[2103] = ~(in[171] | in[139]); 
    assign layer_0[2104] = in[252]; 
    assign layer_0[2105] = in[149] & ~in[9]; 
    assign layer_0[2106] = in[213] | in[182]; 
    assign layer_0[2107] = in[104] ^ in[119]; 
    assign layer_0[2108] = in[183]; 
    assign layer_0[2109] = ~(in[42] | in[51]); 
    assign layer_0[2110] = in[54] ^ in[150]; 
    assign layer_0[2111] = in[93] ^ in[151]; 
    assign layer_0[2112] = in[103]; 
    assign layer_0[2113] = ~(in[85] | in[243]); 
    assign layer_0[2114] = ~(in[118] ^ in[147]); 
    assign layer_0[2115] = in[103] ^ in[211]; 
    assign layer_0[2116] = ~in[229]; 
    assign layer_0[2117] = in[163] | in[145]; 
    assign layer_0[2118] = in[183] & ~in[79]; 
    assign layer_0[2119] = in[79]; 
    assign layer_0[2120] = ~(in[235] ^ in[206]); 
    assign layer_0[2121] = in[131] & ~in[183]; 
    assign layer_0[2122] = in[244] ^ in[247]; 
    assign layer_0[2123] = in[200] | in[131]; 
    assign layer_0[2124] = in[236] | in[148]; 
    assign layer_0[2125] = ~(in[54] ^ in[215]); 
    assign layer_0[2126] = in[93] & ~in[43]; 
    assign layer_0[2127] = ~(in[23] | in[211]); 
    assign layer_0[2128] = in[167] ^ in[185]; 
    assign layer_0[2129] = ~(in[135] ^ in[166]); 
    assign layer_0[2130] = in[43] ^ in[75]; 
    assign layer_0[2131] = in[175] | in[207]; 
    assign layer_0[2132] = ~in[87] | (in[87] & in[166]); 
    assign layer_0[2133] = in[170]; 
    assign layer_0[2134] = ~in[28]; 
    assign layer_0[2135] = in[138]; 
    assign layer_0[2136] = ~(in[98] | in[99]); 
    assign layer_0[2137] = in[140]; 
    assign layer_0[2138] = in[68] & ~in[34]; 
    assign layer_0[2139] = ~(in[143] | in[10]); 
    assign layer_0[2140] = in[214] | in[228]; 
    assign layer_0[2141] = in[8]; 
    assign layer_0[2142] = ~(in[184] ^ in[181]); 
    assign layer_0[2143] = in[156] | in[142]; 
    assign layer_0[2144] = in[100] ^ in[114]; 
    assign layer_0[2145] = ~(in[27] | in[242]); 
    assign layer_0[2146] = ~in[196] | (in[196] & in[98]); 
    assign layer_0[2147] = ~(in[38] ^ in[155]); 
    assign layer_0[2148] = in[149] ^ in[146]; 
    assign layer_0[2149] = ~(in[99] ^ in[97]); 
    assign layer_0[2150] = in[82] ^ in[194]; 
    assign layer_0[2151] = ~in[142] | (in[206] & in[142]); 
    assign layer_0[2152] = in[21]; 
    assign layer_0[2153] = ~(in[90] ^ in[137]); 
    assign layer_0[2154] = ~(in[202] ^ in[235]); 
    assign layer_0[2155] = in[107] ^ in[94]; 
    assign layer_0[2156] = ~(in[219] ^ in[188]); 
    assign layer_0[2157] = ~(in[252] ^ in[203]); 
    assign layer_0[2158] = in[169] | in[82]; 
    assign layer_0[2159] = in[170] ^ in[167]; 
    assign layer_0[2160] = in[132] & ~in[249]; 
    assign layer_0[2161] = ~(in[194] | in[221]); 
    assign layer_0[2162] = ~(in[190] ^ in[221]); 
    assign layer_0[2163] = in[228] | in[72]; 
    assign layer_0[2164] = ~(in[141] ^ in[123]); 
    assign layer_0[2165] = in[203] | in[225]; 
    assign layer_0[2166] = in[221]; 
    assign layer_0[2167] = ~(in[211] ^ in[243]); 
    assign layer_0[2168] = ~(in[189] | in[247]); 
    assign layer_0[2169] = ~(in[23] ^ in[221]); 
    assign layer_0[2170] = in[246] & ~in[177]; 
    assign layer_0[2171] = in[150] & ~in[210]; 
    assign layer_0[2172] = in[72] & ~in[151]; 
    assign layer_0[2173] = ~(in[22] ^ in[53]); 
    assign layer_0[2174] = ~(in[45] ^ in[26]); 
    assign layer_0[2175] = ~in[71]; 
    assign layer_0[2176] = ~(in[196] ^ in[198]); 
    assign layer_0[2177] = in[93] ^ in[75]; 
    assign layer_0[2178] = ~(in[233] | in[218]); 
    assign layer_0[2179] = in[139] & ~in[213]; 
    assign layer_0[2180] = in[38] ^ in[195]; 
    assign layer_0[2181] = in[89] ^ in[220]; 
    assign layer_0[2182] = ~(in[87] ^ in[146]); 
    assign layer_0[2183] = ~(in[184] ^ in[149]); 
    assign layer_0[2184] = ~(in[164] ^ in[199]); 
    assign layer_0[2185] = in[113] | in[114]; 
    assign layer_0[2186] = ~in[126] | (in[251] & in[126]); 
    assign layer_0[2187] = in[187] | in[12]; 
    assign layer_0[2188] = in[211] ^ in[5]; 
    assign layer_0[2189] = ~(in[115] ^ in[41]); 
    assign layer_0[2190] = ~in[57] | (in[57] & in[116]); 
    assign layer_0[2191] = in[206] | in[204]; 
    assign layer_0[2192] = ~(in[237] | in[146]); 
    assign layer_0[2193] = in[211] ^ in[181]; 
    assign layer_0[2194] = ~(in[246] ^ in[55]); 
    assign layer_0[2195] = in[126] | in[182]; 
    assign layer_0[2196] = in[166] ^ in[186]; 
    assign layer_0[2197] = in[211] | in[39]; 
    assign layer_0[2198] = in[57] ^ in[55]; 
    assign layer_0[2199] = ~in[90] | (in[40] & in[90]); 
    assign layer_0[2200] = in[137]; 
    assign layer_0[2201] = in[125] | in[252]; 
    assign layer_0[2202] = in[170] ^ in[83]; 
    assign layer_0[2203] = in[187]; 
    assign layer_0[2204] = ~in[135]; 
    assign layer_0[2205] = in[243]; 
    assign layer_0[2206] = in[247] | in[53]; 
    assign layer_0[2207] = in[241] | in[245]; 
    assign layer_0[2208] = in[149]; 
    assign layer_0[2209] = ~in[125] | (in[125] & in[134]); 
    assign layer_0[2210] = ~in[138] | (in[138] & in[195]); 
    assign layer_0[2211] = in[199] ^ in[156]; 
    assign layer_0[2212] = ~(in[146] | in[150]); 
    assign layer_0[2213] = in[204] ^ in[234]; 
    assign layer_0[2214] = in[197] ^ in[44]; 
    assign layer_0[2215] = in[35] | in[60]; 
    assign layer_0[2216] = in[149] | in[153]; 
    assign layer_0[2217] = ~(in[235] | in[106]); 
    assign layer_0[2218] = ~(in[131] | in[180]); 
    assign layer_0[2219] = in[174] ^ in[7]; 
    assign layer_0[2220] = ~in[133] | (in[99] & in[133]); 
    assign layer_0[2221] = ~(in[98] ^ in[85]); 
    assign layer_0[2222] = ~(in[212] | in[5]); 
    assign layer_0[2223] = ~(in[218] | in[220]); 
    assign layer_0[2224] = in[119] ^ in[84]; 
    assign layer_0[2225] = in[86] ^ in[41]; 
    assign layer_0[2226] = ~(in[6] | in[135]); 
    assign layer_0[2227] = in[81] | in[91]; 
    assign layer_0[2228] = ~(in[120] | in[104]); 
    assign layer_0[2229] = in[101] | in[56]; 
    assign layer_0[2230] = in[56] ^ in[25]; 
    assign layer_0[2231] = ~(in[74] ^ in[43]); 
    assign layer_0[2232] = ~(in[109] ^ in[50]); 
    assign layer_0[2233] = ~(in[125] ^ in[121]); 
    assign layer_0[2234] = ~in[232] | (in[232] & in[108]); 
    assign layer_0[2235] = in[106] ^ in[138]; 
    assign layer_0[2236] = ~(in[183] | in[197]); 
    assign layer_0[2237] = ~(in[93] ^ in[91]); 
    assign layer_0[2238] = ~(in[87] ^ in[168]); 
    assign layer_0[2239] = in[179] & ~in[250]; 
    assign layer_0[2240] = ~in[154] | (in[11] & in[154]); 
    assign layer_0[2241] = in[199] & ~in[147]; 
    assign layer_0[2242] = in[141] ^ in[190]; 
    assign layer_0[2243] = in[247] ^ in[93]; 
    assign layer_0[2244] = ~(in[11] ^ in[42]); 
    assign layer_0[2245] = in[183] & ~in[171]; 
    assign layer_0[2246] = in[151] & ~in[184]; 
    assign layer_0[2247] = in[101] & ~in[172]; 
    assign layer_0[2248] = ~(in[36] ^ in[104]); 
    assign layer_0[2249] = ~(in[182] ^ in[185]); 
    assign layer_0[2250] = in[74] ^ in[172]; 
    assign layer_0[2251] = in[156] ^ in[158]; 
    assign layer_0[2252] = ~(in[63] ^ in[114]); 
    assign layer_0[2253] = in[183] & ~in[90]; 
    assign layer_0[2254] = in[241] | in[105]; 
    assign layer_0[2255] = in[154] ^ in[119]; 
    assign layer_0[2256] = ~(in[106] ^ in[108]); 
    assign layer_0[2257] = in[61] & ~in[217]; 
    assign layer_0[2258] = ~in[101] | (in[197] & in[101]); 
    assign layer_0[2259] = in[71] & ~in[46]; 
    assign layer_0[2260] = in[165] ^ in[196]; 
    assign layer_0[2261] = in[154] | in[133]; 
    assign layer_0[2262] = ~(in[84] | in[147]); 
    assign layer_0[2263] = ~(in[56] ^ in[88]); 
    assign layer_0[2264] = in[92]; 
    assign layer_0[2265] = ~in[204]; 
    assign layer_0[2266] = in[83] & ~in[165]; 
    assign layer_0[2267] = in[8]; 
    assign layer_0[2268] = ~(in[220] ^ in[235]); 
    assign layer_0[2269] = ~in[71] | (in[74] & in[71]); 
    assign layer_0[2270] = ~(in[152] ^ in[121]); 
    assign layer_0[2271] = ~(in[113] ^ in[137]); 
    assign layer_0[2272] = in[179] & ~in[220]; 
    assign layer_0[2273] = in[194]; 
    assign layer_0[2274] = in[198] & ~in[243]; 
    assign layer_0[2275] = ~(in[71] ^ in[41]); 
    assign layer_0[2276] = ~(in[234] | in[212]); 
    assign layer_0[2277] = ~(in[155] | in[53]); 
    assign layer_0[2278] = ~(in[210] | in[143]); 
    assign layer_0[2279] = ~(in[45] ^ in[79]); 
    assign layer_0[2280] = in[147] ^ in[43]; 
    assign layer_0[2281] = in[242] | in[243]; 
    assign layer_0[2282] = ~(in[155] ^ in[142]); 
    assign layer_0[2283] = ~(in[227] | in[23]); 
    assign layer_0[2284] = in[27] & ~in[136]; 
    assign layer_0[2285] = ~(in[118] ^ in[70]); 
    assign layer_0[2286] = ~in[229]; 
    assign layer_0[2287] = ~(in[235] | in[204]); 
    assign layer_0[2288] = in[101] ^ in[35]; 
    assign layer_0[2289] = in[151] & ~in[68]; 
    assign layer_0[2290] = in[39] ^ in[37]; 
    assign layer_0[2291] = in[69] & in[57]; 
    assign layer_0[2292] = ~(in[201] | in[39]); 
    assign layer_0[2293] = in[242] | in[218]; 
    assign layer_0[2294] = in[178] | in[230]; 
    assign layer_0[2295] = ~(in[11] | in[9]); 
    assign layer_0[2296] = ~in[152] | (in[152] & in[171]); 
    assign layer_0[2297] = in[196] | in[178]; 
    assign layer_0[2298] = ~(in[165] ^ in[183]); 
    assign layer_0[2299] = in[87] ^ in[57]; 
    assign layer_0[2300] = ~in[118] | (in[118] & in[10]); 
    assign layer_0[2301] = in[233] ^ in[216]; 
    assign layer_0[2302] = ~(in[116] ^ in[102]); 
    assign layer_0[2303] = in[84] & in[117]; 
    assign layer_0[2304] = ~(in[87] ^ in[67]); 
    assign layer_0[2305] = ~(in[74] ^ in[122]); 
    assign layer_0[2306] = in[149]; 
    assign layer_0[2307] = ~(in[63] ^ in[75]); 
    assign layer_0[2308] = ~(in[159] | in[218]); 
    assign layer_0[2309] = ~(in[53] ^ in[107]); 
    assign layer_0[2310] = in[143] | in[36]; 
    assign layer_0[2311] = in[49] | in[141]; 
    assign layer_0[2312] = in[12] | in[5]; 
    assign layer_0[2313] = in[68] & ~in[240]; 
    assign layer_0[2314] = ~(in[217] ^ in[249]); 
    assign layer_0[2315] = ~(in[200] ^ in[247]); 
    assign layer_0[2316] = in[139] | in[157]; 
    assign layer_0[2317] = in[211] ^ in[151]; 
    assign layer_0[2318] = in[70] | in[241]; 
    assign layer_0[2319] = in[198] ^ in[115]; 
    assign layer_0[2320] = ~(in[93] ^ in[155]); 
    assign layer_0[2321] = ~in[74]; 
    assign layer_0[2322] = ~(in[37] | in[24]); 
    assign layer_0[2323] = ~in[87]; 
    assign layer_0[2324] = in[204] ^ in[201]; 
    assign layer_0[2325] = ~in[184] | (in[184] & in[251]); 
    assign layer_0[2326] = ~(in[46] | in[143]); 
    assign layer_0[2327] = ~(in[110] | in[109]); 
    assign layer_0[2328] = in[132] & ~in[103]; 
    assign layer_0[2329] = in[237] ^ in[206]; 
    assign layer_0[2330] = ~(in[127] ^ in[22]); 
    assign layer_0[2331] = ~(in[121] ^ in[171]); 
    assign layer_0[2332] = ~(in[95] ^ in[63]); 
    assign layer_0[2333] = ~(in[164] | in[146]); 
    assign layer_0[2334] = in[186] | in[218]; 
    assign layer_0[2335] = ~(in[65] | in[152]); 
    assign layer_0[2336] = ~(in[57] ^ in[25]); 
    assign layer_0[2337] = ~(in[196] ^ in[203]); 
    assign layer_0[2338] = in[214]; 
    assign layer_0[2339] = in[214] ^ in[245]; 
    assign layer_0[2340] = ~(in[25] ^ in[55]); 
    assign layer_0[2341] = ~in[52] | (in[52] & in[187]); 
    assign layer_0[2342] = in[103] | in[235]; 
    assign layer_0[2343] = in[78] ^ in[76]; 
    assign layer_0[2344] = in[44] | in[59]; 
    assign layer_0[2345] = in[210] ^ in[100]; 
    assign layer_0[2346] = in[169]; 
    assign layer_0[2347] = in[179] ^ in[181]; 
    assign layer_0[2348] = in[25] & ~in[88]; 
    assign layer_0[2349] = ~(in[143] ^ in[205]); 
    assign layer_0[2350] = ~(in[9] ^ in[196]); 
    assign layer_0[2351] = ~(in[69] ^ in[22]); 
    assign layer_0[2352] = ~(in[196] | in[212]); 
    assign layer_0[2353] = in[139] ^ in[134]; 
    assign layer_0[2354] = in[151] | in[133]; 
    assign layer_0[2355] = in[211] | in[166]; 
    assign layer_0[2356] = ~(in[91] ^ in[109]); 
    assign layer_0[2357] = ~(in[5] ^ in[6]); 
    assign layer_0[2358] = in[181] ^ in[229]; 
    assign layer_0[2359] = ~in[41] | (in[12] & in[41]); 
    assign layer_0[2360] = ~(in[4] | in[27]); 
    assign layer_0[2361] = ~(in[196] ^ in[136]); 
    assign layer_0[2362] = ~in[55]; 
    assign layer_0[2363] = in[196] ^ in[205]; 
    assign layer_0[2364] = ~(in[35] | in[236]); 
    assign layer_0[2365] = ~(in[65] ^ in[168]); 
    assign layer_0[2366] = ~in[136] | (in[165] & in[136]); 
    assign layer_0[2367] = ~in[135] | (in[135] & in[140]); 
    assign layer_0[2368] = in[166] ^ in[184]; 
    assign layer_0[2369] = ~(in[247] | in[110]); 
    assign layer_0[2370] = ~(in[221] ^ in[12]); 
    assign layer_0[2371] = ~in[212]; 
    assign layer_0[2372] = ~(in[185] ^ in[232]); 
    assign layer_0[2373] = ~(in[158] | in[198]); 
    assign layer_0[2374] = ~(in[66] ^ in[38]); 
    assign layer_0[2375] = in[242] | in[242]; 
    assign layer_0[2376] = in[21]; 
    assign layer_0[2377] = ~(in[200] | in[233]); 
    assign layer_0[2378] = in[57] & ~in[171]; 
    assign layer_0[2379] = ~(in[149] | in[151]); 
    assign layer_0[2380] = ~in[119] | (in[162] & in[119]); 
    assign layer_0[2381] = ~(in[150] | in[119]); 
    assign layer_0[2382] = in[94] | in[141]; 
    assign layer_0[2383] = in[109]; 
    assign layer_0[2384] = in[131] ^ in[148]; 
    assign layer_0[2385] = ~in[195] | (in[195] & in[117]); 
    assign layer_0[2386] = ~(in[242] | in[85]); 
    assign layer_0[2387] = in[8] | in[6]; 
    assign layer_0[2388] = ~(in[197] ^ in[162]); 
    assign layer_0[2389] = ~(in[72] ^ in[40]); 
    assign layer_0[2390] = in[131] | in[54]; 
    assign layer_0[2391] = in[215] & ~in[107]; 
    assign layer_0[2392] = ~(in[73] | in[34]); 
    assign layer_0[2393] = in[103] & ~in[6]; 
    assign layer_0[2394] = ~in[108]; 
    assign layer_0[2395] = in[21] & ~in[99]; 
    assign layer_0[2396] = in[24] & ~in[69]; 
    assign layer_0[2397] = in[152]; 
    assign layer_0[2398] = ~in[158]; 
    assign layer_0[2399] = ~in[102] | (in[204] & in[102]); 
    assign layer_0[2400] = in[83] ^ in[165]; 
    assign layer_0[2401] = in[74] | in[210]; 
    assign layer_0[2402] = in[247] | in[39]; 
    assign layer_0[2403] = in[58] ^ in[233]; 
    assign layer_0[2404] = ~in[126] | (in[74] & in[126]); 
    assign layer_0[2405] = ~(in[174] | in[193]); 
    assign layer_0[2406] = ~(in[44] ^ in[106]); 
    assign layer_0[2407] = in[247] & ~in[197]; 
    assign layer_0[2408] = ~in[140] | (in[216] & in[140]); 
    assign layer_0[2409] = ~(in[102] ^ in[140]); 
    assign layer_0[2410] = ~in[88]; 
    assign layer_0[2411] = ~(in[63] | in[100]); 
    assign layer_0[2412] = ~(in[58] ^ in[90]); 
    assign layer_0[2413] = ~in[58] | (in[24] & in[58]); 
    assign layer_0[2414] = in[84] ^ in[71]; 
    assign layer_0[2415] = in[83] & ~in[144]; 
    assign layer_0[2416] = ~(in[155] | in[185]); 
    assign layer_0[2417] = in[169]; 
    assign layer_0[2418] = in[149] & ~in[170]; 
    assign layer_0[2419] = ~(in[155] | in[171]); 
    assign layer_0[2420] = ~in[88]; 
    assign layer_0[2421] = ~(in[151] ^ in[227]); 
    assign layer_0[2422] = in[106] | in[124]; 
    assign layer_0[2423] = in[119] | in[135]; 
    assign layer_0[2424] = ~(in[181] ^ in[202]); 
    assign layer_0[2425] = ~(in[122] | in[140]); 
    assign layer_0[2426] = ~in[196] | (in[196] & in[210]); 
    assign layer_0[2427] = ~(in[113] ^ in[100]); 
    assign layer_0[2428] = in[119]; 
    assign layer_0[2429] = in[125] | in[139]; 
    assign layer_0[2430] = ~in[101] | (in[104] & in[101]); 
    assign layer_0[2431] = ~(in[151] ^ in[121]); 
    assign layer_0[2432] = ~(in[149] | in[162]); 
    assign layer_0[2433] = ~in[120]; 
    assign layer_0[2434] = in[109] | in[181]; 
    assign layer_0[2435] = in[10] | in[30]; 
    assign layer_0[2436] = in[218] & ~in[124]; 
    assign layer_0[2437] = in[116] ^ in[130]; 
    assign layer_0[2438] = ~(in[186] | in[203]); 
    assign layer_0[2439] = ~(in[199] | in[135]); 
    assign layer_0[2440] = in[148] | in[115]; 
    assign layer_0[2441] = in[177] | in[148]; 
    assign layer_0[2442] = in[72] & ~in[27]; 
    assign layer_0[2443] = in[161] | in[193]; 
    assign layer_0[2444] = ~(in[23] | in[184]); 
    assign layer_0[2445] = ~(in[152] | in[78]); 
    assign layer_0[2446] = ~(in[27] ^ in[107]); 
    assign layer_0[2447] = in[182] | in[196]; 
    assign layer_0[2448] = in[216]; 
    assign layer_0[2449] = ~(in[29] ^ in[63]); 
    assign layer_0[2450] = in[248] ^ in[216]; 
    assign layer_0[2451] = in[229] | in[177]; 
    assign layer_0[2452] = ~in[50]; 
    assign layer_0[2453] = in[39] ^ in[69]; 
    assign layer_0[2454] = ~(in[169] ^ in[172]); 
    assign layer_0[2455] = in[36]; 
    assign layer_0[2456] = ~in[189]; 
    assign layer_0[2457] = ~(in[75] | in[147]); 
    assign layer_0[2458] = in[68] ^ in[37]; 
    assign layer_0[2459] = in[233] ^ in[197]; 
    assign layer_0[2460] = in[52] | in[194]; 
    assign layer_0[2461] = ~(in[142] | in[132]); 
    assign layer_0[2462] = ~in[104] | (in[195] & in[104]); 
    assign layer_0[2463] = in[121]; 
    assign layer_0[2464] = ~in[119]; 
    assign layer_0[2465] = ~in[138] | (in[9] & in[138]); 
    assign layer_0[2466] = ~(in[121] ^ in[146]); 
    assign layer_0[2467] = in[73] ^ in[70]; 
    assign layer_0[2468] = in[88] | in[184]; 
    assign layer_0[2469] = ~(in[30] | in[115]); 
    assign layer_0[2470] = in[8] ^ in[188]; 
    assign layer_0[2471] = ~(in[250] | in[135]); 
    assign layer_0[2472] = ~(in[169] | in[171]); 
    assign layer_0[2473] = ~(in[141] ^ in[108]); 
    assign layer_0[2474] = ~(in[60] | in[53]); 
    assign layer_0[2475] = in[71] ^ in[213]; 
    assign layer_0[2476] = ~in[104] | (in[104] & in[88]); 
    assign layer_0[2477] = ~(in[118] | in[212]); 
    assign layer_0[2478] = ~in[108] | (in[108] & in[89]); 
    assign layer_0[2479] = ~in[101] | (in[101] & in[211]); 
    assign layer_0[2480] = in[63] ^ in[100]; 
    assign layer_0[2481] = in[122] ^ in[124]; 
    assign layer_0[2482] = in[108] ^ in[140]; 
    assign layer_0[2483] = ~in[55] | (in[21] & in[55]); 
    assign layer_0[2484] = ~(in[104] ^ in[136]); 
    assign layer_0[2485] = in[228] & ~in[187]; 
    assign layer_0[2486] = ~(in[107] | in[125]); 
    assign layer_0[2487] = ~(in[195] ^ in[100]); 
    assign layer_0[2488] = in[203]; 
    assign layer_0[2489] = ~(in[139] ^ in[23]); 
    assign layer_0[2490] = in[136]; 
    assign layer_0[2491] = in[183] ^ in[232]; 
    assign layer_0[2492] = ~in[179]; 
    assign layer_0[2493] = in[137] ^ in[105]; 
    assign layer_0[2494] = in[34] | in[186]; 
    assign layer_0[2495] = in[19]; 
    assign layer_0[2496] = ~(in[205] | in[26]); 
    assign layer_0[2497] = in[10] ^ in[29]; 
    assign layer_0[2498] = ~in[242]; 
    assign layer_0[2499] = in[11] | in[242]; 
    assign layer_0[2500] = ~(in[6] ^ in[139]); 
    assign layer_0[2501] = ~(in[158] ^ in[141]); 
    assign layer_0[2502] = ~(in[30] | in[52]); 
    assign layer_0[2503] = in[213] ^ in[243]; 
    assign layer_0[2504] = ~in[235]; 
    assign layer_0[2505] = ~(in[45] | in[79]); 
    assign layer_0[2506] = ~(in[175] | in[203]); 
    assign layer_0[2507] = in[215] & ~in[55]; 
    assign layer_0[2508] = in[181] ^ in[139]; 
    assign layer_0[2509] = in[78] | in[199]; 
    assign layer_0[2510] = ~(in[169] | in[138]); 
    assign layer_0[2511] = in[40] ^ in[122]; 
    assign layer_0[2512] = in[50] | in[81]; 
    assign layer_0[2513] = in[229] | in[25]; 
    assign layer_0[2514] = ~(in[71] | in[40]); 
    assign layer_0[2515] = in[204]; 
    assign layer_0[2516] = in[136]; 
    assign layer_0[2517] = in[103] ^ in[89]; 
    assign layer_0[2518] = in[220] ^ in[250]; 
    assign layer_0[2519] = ~(in[75] ^ in[155]); 
    assign layer_0[2520] = in[52] | in[187]; 
    assign layer_0[2521] = in[88] | in[92]; 
    assign layer_0[2522] = in[248] | in[87]; 
    assign layer_0[2523] = in[150] ^ in[151]; 
    assign layer_0[2524] = in[163] | in[148]; 
    assign layer_0[2525] = ~(in[103] | in[29]); 
    assign layer_0[2526] = ~(in[56] | in[237]); 
    assign layer_0[2527] = ~(in[102] ^ in[88]); 
    assign layer_0[2528] = in[99] | in[170]; 
    assign layer_0[2529] = in[140] & ~in[200]; 
    assign layer_0[2530] = ~in[245]; 
    assign layer_0[2531] = in[55] ^ in[24]; 
    assign layer_0[2532] = in[68] | in[42]; 
    assign layer_0[2533] = in[129] | in[34]; 
    assign layer_0[2534] = ~(in[154] ^ in[21]); 
    assign layer_0[2535] = ~(in[146] | in[242]); 
    assign layer_0[2536] = in[131] & ~in[153]; 
    assign layer_0[2537] = in[133] & ~in[35]; 
    assign layer_0[2538] = in[79] & ~in[19]; 
    assign layer_0[2539] = in[118] ^ in[126]; 
    assign layer_0[2540] = ~in[141]; 
    assign layer_0[2541] = in[79] | in[248]; 
    assign layer_0[2542] = ~(in[120] & in[123]); 
    assign layer_0[2543] = in[53] & ~in[202]; 
    assign layer_0[2544] = ~(in[162] & in[162]); 
    assign layer_0[2545] = in[50] | in[26]; 
    assign layer_0[2546] = ~(in[103] | in[72]); 
    assign layer_0[2547] = in[166] & ~in[245]; 
    assign layer_0[2548] = in[210] ^ in[72]; 
    assign layer_0[2549] = in[118] ^ in[52]; 
    assign layer_0[2550] = in[122] & ~in[9]; 
    assign layer_0[2551] = in[61] ^ in[78]; 
    assign layer_0[2552] = in[49] | in[84]; 
    assign layer_0[2553] = in[118] | in[131]; 
    assign layer_0[2554] = in[163] | in[130]; 
    assign layer_0[2555] = ~(in[142] | in[143]); 
    assign layer_0[2556] = ~(in[218] | in[52]); 
    assign layer_0[2557] = in[247] ^ in[215]; 
    assign layer_0[2558] = in[231] ^ in[216]; 
    assign layer_0[2559] = ~(in[140] | in[187]); 
    // Layer 1 ============================================================
    assign out[0] = ~layer_0[1447] | (layer_0[1447] & layer_0[681]); 
    assign out[1] = layer_0[1911] & ~layer_0[1141]; 
    assign out[2] = ~(layer_0[1215] | layer_0[758]); 
    assign out[3] = ~(layer_0[1629] ^ layer_0[1]); 
    assign out[4] = layer_0[278]; 
    assign out[5] = layer_0[2339]; 
    assign out[6] = ~layer_0[2074]; 
    assign out[7] = ~layer_0[1810] | (layer_0[1810] & layer_0[1555]); 
    assign out[8] = layer_0[1108] & ~layer_0[2512]; 
    assign out[9] = layer_0[1558] & ~layer_0[2164]; 
    assign out[10] = layer_0[312] | layer_0[1983]; 
    assign out[11] = ~(layer_0[684] ^ layer_0[957]); 
    assign out[12] = layer_0[1021]; 
    assign out[13] = layer_0[1918] & layer_0[661]; 
    assign out[14] = layer_0[833] ^ layer_0[843]; 
    assign out[15] = layer_0[1660] ^ layer_0[451]; 
    assign out[16] = ~layer_0[2053]; 
    assign out[17] = layer_0[1895] ^ layer_0[679]; 
    assign out[18] = ~layer_0[1465]; 
    assign out[19] = layer_0[364] ^ layer_0[790]; 
    assign out[20] = layer_0[1143] & ~layer_0[1474]; 
    assign out[21] = layer_0[1906] & layer_0[991]; 
    assign out[22] = layer_0[1571]; 
    assign out[23] = ~(layer_0[2260] ^ layer_0[2440]); 
    assign out[24] = ~(layer_0[1903] | layer_0[878]); 
    assign out[25] = ~(layer_0[1238] ^ layer_0[688]); 
    assign out[26] = ~layer_0[1585]; 
    assign out[27] = ~layer_0[48]; 
    assign out[28] = ~layer_0[773]; 
    assign out[29] = ~layer_0[2235]; 
    assign out[30] = ~(layer_0[159] ^ layer_0[1587]); 
    assign out[31] = layer_0[2272]; 
    assign out[32] = layer_0[2018]; 
    assign out[33] = layer_0[1849] | layer_0[817]; 
    assign out[34] = layer_0[3] & ~layer_0[2196]; 
    assign out[35] = ~(layer_0[1395] & layer_0[1039]); 
    assign out[36] = ~layer_0[1003]; 
    assign out[37] = ~layer_0[1970]; 
    assign out[38] = layer_0[1849] & layer_0[561]; 
    assign out[39] = layer_0[1694]; 
    assign out[40] = layer_0[2169] ^ layer_0[740]; 
    assign out[41] = layer_0[2153] & ~layer_0[607]; 
    assign out[42] = layer_0[2043] ^ layer_0[2223]; 
    assign out[43] = ~layer_0[209]; 
    assign out[44] = ~layer_0[1589]; 
    assign out[45] = ~(layer_0[1051] | layer_0[390]); 
    assign out[46] = ~layer_0[1183] | (layer_0[260] & layer_0[1183]); 
    assign out[47] = layer_0[1233] ^ layer_0[1809]; 
    assign out[48] = layer_0[1319] & ~layer_0[6]; 
    assign out[49] = layer_0[1849] & layer_0[1041]; 
    assign out[50] = layer_0[1766]; 
    assign out[51] = ~(layer_0[1836] | layer_0[875]); 
    assign out[52] = layer_0[2155] & layer_0[2440]; 
    assign out[53] = layer_0[1414] & ~layer_0[899]; 
    assign out[54] = layer_0[276] & ~layer_0[1776]; 
    assign out[55] = layer_0[3] & ~layer_0[1111]; 
    assign out[56] = layer_0[789] ^ layer_0[2002]; 
    assign out[57] = layer_0[946] & ~layer_0[760]; 
    assign out[58] = ~layer_0[2255]; 
    assign out[59] = ~(layer_0[1131] ^ layer_0[1386]); 
    assign out[60] = layer_0[1390]; 
    assign out[61] = layer_0[461]; 
    assign out[62] = ~(layer_0[1988] ^ layer_0[1572]); 
    assign out[63] = ~layer_0[1436]; 
    assign out[64] = layer_0[0] & ~layer_0[1632]; 
    assign out[65] = layer_0[2270] & layer_0[661]; 
    assign out[66] = ~(layer_0[816] ^ layer_0[1653]); 
    assign out[67] = ~(layer_0[764] | layer_0[1886]); 
    assign out[68] = ~layer_0[2518]; 
    assign out[69] = layer_0[2172]; 
    assign out[70] = ~layer_0[1810]; 
    assign out[71] = layer_0[871] & ~layer_0[564]; 
    assign out[72] = ~(layer_0[1417] ^ layer_0[715]); 
    assign out[73] = ~layer_0[640]; 
    assign out[74] = ~(layer_0[339] ^ layer_0[939]); 
    assign out[75] = ~layer_0[189]; 
    assign out[76] = ~layer_0[1448]; 
    assign out[77] = layer_0[134] & layer_0[1740]; 
    assign out[78] = ~(layer_0[2453] | layer_0[436]); 
    assign out[79] = layer_0[1532] ^ layer_0[1382]; 
    assign out[80] = layer_0[335] & layer_0[205]; 
    assign out[81] = ~layer_0[145] | (layer_0[1147] & layer_0[145]); 
    assign out[82] = layer_0[783] & layer_0[1752]; 
    assign out[83] = layer_0[2510]; 
    assign out[84] = ~layer_0[839] | (layer_0[1416] & layer_0[839]); 
    assign out[85] = layer_0[1068] ^ layer_0[2066]; 
    assign out[86] = ~layer_0[2555] | (layer_0[200] & layer_0[2555]); 
    assign out[87] = layer_0[77] & ~layer_0[740]; 
    assign out[88] = layer_0[2173] & ~layer_0[2307]; 
    assign out[89] = layer_0[2129]; 
    assign out[90] = ~(layer_0[892] | layer_0[420]); 
    assign out[91] = ~layer_0[1773] | (layer_0[1372] & layer_0[1773]); 
    assign out[92] = layer_0[1547] & ~layer_0[1721]; 
    assign out[93] = layer_0[1520] ^ layer_0[831]; 
    assign out[94] = layer_0[2190] ^ layer_0[1572]; 
    assign out[95] = layer_0[1391] & ~layer_0[990]; 
    assign out[96] = ~layer_0[20] | (layer_0[20] & layer_0[1469]); 
    assign out[97] = ~layer_0[1061]; 
    assign out[98] = layer_0[1052]; 
    assign out[99] = ~layer_0[1603]; 
    assign out[100] = ~(layer_0[1146] ^ layer_0[1258]); 
    assign out[101] = layer_0[938] & layer_0[1155]; 
    assign out[102] = layer_0[1149] ^ layer_0[1481]; 
    assign out[103] = layer_0[1000] & ~layer_0[726]; 
    assign out[104] = ~(layer_0[589] ^ layer_0[2186]); 
    assign out[105] = layer_0[1446]; 
    assign out[106] = layer_0[2182] & layer_0[1918]; 
    assign out[107] = layer_0[1108] & ~layer_0[1706]; 
    assign out[108] = ~layer_0[1164]; 
    assign out[109] = ~(layer_0[9] | layer_0[1115]); 
    assign out[110] = layer_0[807] & ~layer_0[2435]; 
    assign out[111] = layer_0[2384]; 
    assign out[112] = layer_0[1901]; 
    assign out[113] = ~(layer_0[162] & layer_0[273]); 
    assign out[114] = layer_0[853] ^ layer_0[319]; 
    assign out[115] = layer_0[857] & ~layer_0[2290]; 
    assign out[116] = layer_0[166] & ~layer_0[1234]; 
    assign out[117] = layer_0[1696] ^ layer_0[403]; 
    assign out[118] = layer_0[2059] & ~layer_0[356]; 
    assign out[119] = layer_0[24] & ~layer_0[1312]; 
    assign out[120] = ~(layer_0[1894] | layer_0[1794]); 
    assign out[121] = layer_0[889]; 
    assign out[122] = ~(layer_0[1565] & layer_0[2327]); 
    assign out[123] = ~(layer_0[2219] ^ layer_0[145]); 
    assign out[124] = ~(layer_0[2489] ^ layer_0[1635]); 
    assign out[125] = ~(layer_0[2484] ^ layer_0[2063]); 
    assign out[126] = layer_0[2297] & layer_0[1618]; 
    assign out[127] = ~layer_0[1465]; 
    assign out[128] = ~layer_0[2235] | (layer_0[2235] & layer_0[1305]); 
    assign out[129] = layer_0[1910]; 
    assign out[130] = ~layer_0[2508]; 
    assign out[131] = ~(layer_0[2266] ^ layer_0[1116]); 
    assign out[132] = ~layer_0[1729]; 
    assign out[133] = layer_0[803] & ~layer_0[863]; 
    assign out[134] = layer_0[705] ^ layer_0[1738]; 
    assign out[135] = ~(layer_0[413] & layer_0[65]); 
    assign out[136] = layer_0[2238]; 
    assign out[137] = layer_0[335] ^ layer_0[2308]; 
    assign out[138] = layer_0[592] & ~layer_0[1153]; 
    assign out[139] = ~layer_0[1831]; 
    assign out[140] = layer_0[1578] ^ layer_0[2535]; 
    assign out[141] = layer_0[1709] ^ layer_0[1294]; 
    assign out[142] = layer_0[276]; 
    assign out[143] = ~layer_0[73]; 
    assign out[144] = ~(layer_0[1153] | layer_0[2158]); 
    assign out[145] = layer_0[264]; 
    assign out[146] = layer_0[2268] & ~layer_0[496]; 
    assign out[147] = ~layer_0[15]; 
    assign out[148] = layer_0[893] & ~layer_0[1641]; 
    assign out[149] = layer_0[372] & ~layer_0[2056]; 
    assign out[150] = layer_0[1143] & ~layer_0[118]; 
    assign out[151] = ~(layer_0[1213] & layer_0[1742]); 
    assign out[152] = ~(layer_0[1052] ^ layer_0[1752]); 
    assign out[153] = layer_0[296]; 
    assign out[154] = layer_0[614] & layer_0[2270]; 
    assign out[155] = ~(layer_0[2493] | layer_0[1200]); 
    assign out[156] = layer_0[1912]; 
    assign out[157] = layer_0[1139] & ~layer_0[1215]; 
    assign out[158] = layer_0[1567]; 
    assign out[159] = ~(layer_0[1431] ^ layer_0[59]); 
    assign out[160] = ~layer_0[345]; 
    assign out[161] = layer_0[176] & layer_0[609]; 
    assign out[162] = layer_0[1532] ^ layer_0[629]; 
    assign out[163] = ~layer_0[2064]; 
    assign out[164] = ~(layer_0[1798] ^ layer_0[1409]); 
    assign out[165] = layer_0[2103] ^ layer_0[1211]; 
    assign out[166] = layer_0[1967] ^ layer_0[2120]; 
    assign out[167] = layer_0[1331] | layer_0[1851]; 
    assign out[168] = ~(layer_0[543] ^ layer_0[2268]); 
    assign out[169] = ~(layer_0[1801] | layer_0[1615]); 
    assign out[170] = ~(layer_0[2453] | layer_0[2235]); 
    assign out[171] = ~(layer_0[1734] ^ layer_0[502]); 
    assign out[172] = layer_0[139] | layer_0[588]; 
    assign out[173] = ~(layer_0[648] | layer_0[1296]); 
    assign out[174] = layer_0[996] ^ layer_0[1175]; 
    assign out[175] = ~(layer_0[1189] ^ layer_0[2425]); 
    assign out[176] = ~(layer_0[1324] & layer_0[713]); 
    assign out[177] = layer_0[1541]; 
    assign out[178] = layer_0[304] ^ layer_0[1356]; 
    assign out[179] = layer_0[457] ^ layer_0[1595]; 
    assign out[180] = ~(layer_0[1894] | layer_0[1193]); 
    assign out[181] = ~(layer_0[1654] | layer_0[2128]); 
    assign out[182] = layer_0[1989]; 
    assign out[183] = layer_0[2120]; 
    assign out[184] = ~(layer_0[515] ^ layer_0[1777]); 
    assign out[185] = ~layer_0[381] | (layer_0[1500] & layer_0[381]); 
    assign out[186] = layer_0[433] & ~layer_0[701]; 
    assign out[187] = layer_0[1333] & layer_0[541]; 
    assign out[188] = ~(layer_0[151] & layer_0[2176]); 
    assign out[189] = layer_0[1974] ^ layer_0[1087]; 
    assign out[190] = ~layer_0[1903] | (layer_0[1903] & layer_0[1710]); 
    assign out[191] = layer_0[942]; 
    assign out[192] = ~layer_0[1723]; 
    assign out[193] = ~layer_0[1292]; 
    assign out[194] = layer_0[989] ^ layer_0[811]; 
    assign out[195] = layer_0[1664] ^ layer_0[2095]; 
    assign out[196] = layer_0[1710]; 
    assign out[197] = ~(layer_0[351] ^ layer_0[2468]); 
    assign out[198] = ~layer_0[2540] | (layer_0[2540] & layer_0[1218]); 
    assign out[199] = ~layer_0[976]; 
    assign out[200] = layer_0[1109] ^ layer_0[1855]; 
    assign out[201] = ~layer_0[714]; 
    assign out[202] = ~(layer_0[132] ^ layer_0[1255]); 
    assign out[203] = layer_0[1627]; 
    assign out[204] = ~(layer_0[2265] ^ layer_0[575]); 
    assign out[205] = layer_0[502] & ~layer_0[1938]; 
    assign out[206] = ~(layer_0[1902] ^ layer_0[2102]); 
    assign out[207] = ~layer_0[1777]; 
    assign out[208] = layer_0[1237]; 
    assign out[209] = ~(layer_0[60] | layer_0[209]); 
    assign out[210] = layer_0[2335] & ~layer_0[898]; 
    assign out[211] = layer_0[592]; 
    assign out[212] = layer_0[2477] ^ layer_0[2034]; 
    assign out[213] = layer_0[2425] & ~layer_0[964]; 
    assign out[214] = ~(layer_0[15] ^ layer_0[102]); 
    assign out[215] = ~(layer_0[600] ^ layer_0[457]); 
    assign out[216] = ~layer_0[162]; 
    assign out[217] = layer_0[2029] & ~layer_0[1119]; 
    assign out[218] = ~layer_0[839] | (layer_0[839] & layer_0[997]); 
    assign out[219] = ~layer_0[1153]; 
    assign out[220] = ~(layer_0[2255] | layer_0[270]); 
    assign out[221] = layer_0[446]; 
    assign out[222] = ~(layer_0[299] ^ layer_0[1396]); 
    assign out[223] = layer_0[1297] ^ layer_0[1922]; 
    assign out[224] = ~(layer_0[283] | layer_0[684]); 
    assign out[225] = ~layer_0[272] | (layer_0[1021] & layer_0[272]); 
    assign out[226] = ~layer_0[2244] | (layer_0[511] & layer_0[2244]); 
    assign out[227] = ~(layer_0[914] ^ layer_0[2142]); 
    assign out[228] = ~layer_0[277]; 
    assign out[229] = ~(layer_0[401] ^ layer_0[846]); 
    assign out[230] = layer_0[1413] | layer_0[1517]; 
    assign out[231] = layer_0[1569]; 
    assign out[232] = ~layer_0[2255]; 
    assign out[233] = layer_0[1977] & ~layer_0[2428]; 
    assign out[234] = ~(layer_0[457] ^ layer_0[1435]); 
    assign out[235] = layer_0[545] & layer_0[1775]; 
    assign out[236] = layer_0[1633] ^ layer_0[1534]; 
    assign out[237] = layer_0[973]; 
    assign out[238] = layer_0[858] & ~layer_0[78]; 
    assign out[239] = ~(layer_0[301] ^ layer_0[382]); 
    assign out[240] = ~(layer_0[187] ^ layer_0[846]); 
    assign out[241] = layer_0[2086]; 
    assign out[242] = ~(layer_0[1763] | layer_0[1845]); 
    assign out[243] = layer_0[2287] ^ layer_0[40]; 
    assign out[244] = ~layer_0[434]; 
    assign out[245] = layer_0[1850] & ~layer_0[1608]; 
    assign out[246] = layer_0[2071] & ~layer_0[839]; 
    assign out[247] = layer_0[809]; 
    assign out[248] = ~layer_0[1406]; 
    assign out[249] = layer_0[857]; 
    assign out[250] = ~layer_0[1124]; 
    assign out[251] = ~layer_0[2209] | (layer_0[2209] & layer_0[890]); 
    assign out[252] = layer_0[1059] & layer_0[1208]; 
    assign out[253] = ~(layer_0[1888] | layer_0[1483]); 
    assign out[254] = layer_0[569] ^ layer_0[538]; 
    assign out[255] = ~layer_0[2531]; 
    assign out[256] = ~(layer_0[562] & layer_0[2110]); 
    assign out[257] = ~(layer_0[1122] | layer_0[1778]); 
    assign out[258] = ~layer_0[200]; 
    assign out[259] = ~(layer_0[82] | layer_0[1275]); 
    assign out[260] = ~layer_0[1009] | (layer_0[897] & layer_0[1009]); 
    assign out[261] = ~(layer_0[2154] ^ layer_0[562]); 
    assign out[262] = layer_0[36]; 
    assign out[263] = layer_0[1474] ^ layer_0[2277]; 
    assign out[264] = layer_0[2058] ^ layer_0[93]; 
    assign out[265] = layer_0[2176]; 
    assign out[266] = layer_0[1520] ^ layer_0[1507]; 
    assign out[267] = layer_0[2037] & layer_0[760]; 
    assign out[268] = ~layer_0[1784]; 
    assign out[269] = ~layer_0[1293]; 
    assign out[270] = layer_0[301] ^ layer_0[185]; 
    assign out[271] = ~layer_0[335]; 
    assign out[272] = ~layer_0[1934] | (layer_0[2089] & layer_0[1934]); 
    assign out[273] = ~(layer_0[2525] & layer_0[1020]); 
    assign out[274] = ~(layer_0[832] ^ layer_0[1138]); 
    assign out[275] = ~(layer_0[2440] & layer_0[61]); 
    assign out[276] = ~layer_0[626]; 
    assign out[277] = layer_0[1954] & ~layer_0[1520]; 
    assign out[278] = layer_0[1642]; 
    assign out[279] = layer_0[296] ^ layer_0[1871]; 
    assign out[280] = ~layer_0[93]; 
    assign out[281] = layer_0[710]; 
    assign out[282] = layer_0[107] ^ layer_0[1109]; 
    assign out[283] = ~layer_0[66]; 
    assign out[284] = layer_0[2459]; 
    assign out[285] = layer_0[1791] & layer_0[444]; 
    assign out[286] = layer_0[821]; 
    assign out[287] = layer_0[2534] & ~layer_0[1612]; 
    assign out[288] = layer_0[2302] & ~layer_0[567]; 
    assign out[289] = layer_0[1890]; 
    assign out[290] = layer_0[1204] ^ layer_0[1256]; 
    assign out[291] = layer_0[2292] ^ layer_0[804]; 
    assign out[292] = layer_0[303] & layer_0[2490]; 
    assign out[293] = layer_0[170] ^ layer_0[171]; 
    assign out[294] = layer_0[49] & ~layer_0[844]; 
    assign out[295] = layer_0[597] & ~layer_0[1751]; 
    assign out[296] = ~(layer_0[913] | layer_0[2025]); 
    assign out[297] = ~(layer_0[2244] ^ layer_0[1040]); 
    assign out[298] = layer_0[2166]; 
    assign out[299] = layer_0[338]; 
    assign out[300] = layer_0[1922] & layer_0[199]; 
    assign out[301] = layer_0[369] ^ layer_0[793]; 
    assign out[302] = layer_0[1985]; 
    assign out[303] = ~layer_0[1121]; 
    assign out[304] = ~(layer_0[510] ^ layer_0[2204]); 
    assign out[305] = layer_0[710]; 
    assign out[306] = layer_0[2282] & ~layer_0[1401]; 
    assign out[307] = layer_0[1459] ^ layer_0[1972]; 
    assign out[308] = layer_0[117]; 
    assign out[309] = layer_0[1893] ^ layer_0[422]; 
    assign out[310] = ~(layer_0[1870] | layer_0[1253]); 
    assign out[311] = layer_0[1031]; 
    assign out[312] = layer_0[488] ^ layer_0[2356]; 
    assign out[313] = layer_0[2430] & ~layer_0[543]; 
    assign out[314] = ~(layer_0[1095] ^ layer_0[793]); 
    assign out[315] = layer_0[919] & ~layer_0[440]; 
    assign out[316] = ~layer_0[640] | (layer_0[640] & layer_0[1404]); 
    assign out[317] = layer_0[2208] ^ layer_0[719]; 
    assign out[318] = layer_0[1904] & ~layer_0[2547]; 
    assign out[319] = ~(layer_0[384] ^ layer_0[524]); 
    assign out[320] = layer_0[1614] & layer_0[793]; 
    assign out[321] = ~layer_0[588]; 
    assign out[322] = layer_0[1889]; 
    assign out[323] = ~(layer_0[1590] ^ layer_0[1812]); 
    assign out[324] = ~(layer_0[225] | layer_0[277]); 
    assign out[325] = layer_0[997] ^ layer_0[1632]; 
    assign out[326] = layer_0[1035] & layer_0[6]; 
    assign out[327] = ~(layer_0[1936] | layer_0[462]); 
    assign out[328] = ~layer_0[806]; 
    assign out[329] = layer_0[1544] & ~layer_0[2295]; 
    assign out[330] = layer_0[829] & layer_0[1641]; 
    assign out[331] = ~(layer_0[1729] ^ layer_0[899]); 
    assign out[332] = ~(layer_0[2174] | layer_0[2217]); 
    assign out[333] = ~layer_0[2019]; 
    assign out[334] = ~(layer_0[2228] ^ layer_0[1541]); 
    assign out[335] = layer_0[1213]; 
    assign out[336] = layer_0[556]; 
    assign out[337] = ~(layer_0[1648] ^ layer_0[386]); 
    assign out[338] = ~(layer_0[1322] ^ layer_0[1370]); 
    assign out[339] = layer_0[821]; 
    assign out[340] = ~(layer_0[84] ^ layer_0[1017]); 
    assign out[341] = layer_0[399] ^ layer_0[2027]; 
    assign out[342] = layer_0[1794]; 
    assign out[343] = layer_0[574] ^ layer_0[824]; 
    assign out[344] = ~layer_0[63] | (layer_0[63] & layer_0[1580]); 
    assign out[345] = layer_0[1204] | layer_0[449]; 
    assign out[346] = layer_0[2411] & ~layer_0[635]; 
    assign out[347] = ~(layer_0[721] | layer_0[1409]); 
    assign out[348] = layer_0[497] & ~layer_0[1015]; 
    assign out[349] = ~(layer_0[698] ^ layer_0[1324]); 
    assign out[350] = layer_0[1008]; 
    assign out[351] = layer_0[491]; 
    assign out[352] = ~(layer_0[1233] & layer_0[654]); 
    assign out[353] = ~(layer_0[2441] | layer_0[1037]); 
    assign out[354] = layer_0[500] & layer_0[2544]; 
    assign out[355] = layer_0[1201]; 
    assign out[356] = layer_0[2231] & ~layer_0[1583]; 
    assign out[357] = ~(layer_0[1251] | layer_0[66]); 
    assign out[358] = layer_0[2282] & ~layer_0[1325]; 
    assign out[359] = ~(layer_0[939] | layer_0[1869]); 
    assign out[360] = ~(layer_0[2406] ^ layer_0[1717]); 
    assign out[361] = ~layer_0[1991]; 
    assign out[362] = layer_0[602] & ~layer_0[995]; 
    assign out[363] = layer_0[1506] ^ layer_0[1432]; 
    assign out[364] = layer_0[2188] ^ layer_0[1821]; 
    assign out[365] = ~(layer_0[329] ^ layer_0[1493]); 
    assign out[366] = layer_0[763] & ~layer_0[1705]; 
    assign out[367] = ~(layer_0[2180] ^ layer_0[949]); 
    assign out[368] = layer_0[1968] & ~layer_0[1480]; 
    assign out[369] = ~(layer_0[978] & layer_0[2440]); 
    assign out[370] = layer_0[1779] ^ layer_0[424]; 
    assign out[371] = ~(layer_0[1918] ^ layer_0[186]); 
    assign out[372] = ~(layer_0[1874] | layer_0[511]); 
    assign out[373] = layer_0[616]; 
    assign out[374] = layer_0[1110] & layer_0[821]; 
    assign out[375] = layer_0[453]; 
    assign out[376] = layer_0[1845] ^ layer_0[868]; 
    assign out[377] = ~layer_0[873]; 
    assign out[378] = layer_0[35] & layer_0[265]; 
    assign out[379] = layer_0[1444] ^ layer_0[2381]; 
    assign out[380] = layer_0[1757]; 
    assign out[381] = layer_0[2173] ^ layer_0[1319]; 
    assign out[382] = layer_0[2412]; 
    assign out[383] = layer_0[1505] & layer_0[518]; 
    assign out[384] = ~(layer_0[1975] ^ layer_0[1193]); 
    assign out[385] = ~layer_0[737]; 
    assign out[386] = ~(layer_0[1653] ^ layer_0[783]); 
    assign out[387] = ~(layer_0[1880] ^ layer_0[2432]); 
    assign out[388] = layer_0[2305] & ~layer_0[531]; 
    assign out[389] = ~(layer_0[1657] ^ layer_0[2254]); 
    assign out[390] = ~layer_0[2370]; 
    assign out[391] = layer_0[2227] ^ layer_0[602]; 
    assign out[392] = layer_0[2207] ^ layer_0[465]; 
    assign out[393] = layer_0[561] ^ layer_0[766]; 
    assign out[394] = layer_0[129] & layer_0[1882]; 
    assign out[395] = ~(layer_0[1610] ^ layer_0[1995]); 
    assign out[396] = ~layer_0[1004]; 
    assign out[397] = layer_0[2081] & ~layer_0[2531]; 
    assign out[398] = layer_0[57] | layer_0[1947]; 
    assign out[399] = ~(layer_0[1138] ^ layer_0[2021]); 
    assign out[400] = ~(layer_0[236] ^ layer_0[1043]); 
    assign out[401] = layer_0[983] ^ layer_0[1476]; 
    assign out[402] = layer_0[2511]; 
    assign out[403] = layer_0[2282]; 
    assign out[404] = ~layer_0[2506]; 
    assign out[405] = ~(layer_0[1373] | layer_0[2512]); 
    assign out[406] = layer_0[1327] & layer_0[2212]; 
    assign out[407] = ~(layer_0[2233] | layer_0[1919]); 
    assign out[408] = ~(layer_0[1525] ^ layer_0[1806]); 
    assign out[409] = ~layer_0[2183]; 
    assign out[410] = layer_0[2352] ^ layer_0[747]; 
    assign out[411] = ~layer_0[1869]; 
    assign out[412] = layer_0[2115]; 
    assign out[413] = ~(layer_0[486] ^ layer_0[2216]); 
    assign out[414] = layer_0[1042] & layer_0[1172]; 
    assign out[415] = ~(layer_0[670] & layer_0[1126]); 
    assign out[416] = ~layer_0[1792]; 
    assign out[417] = layer_0[1519]; 
    assign out[418] = layer_0[2381] & layer_0[215]; 
    assign out[419] = layer_0[1374] | layer_0[1889]; 
    assign out[420] = ~(layer_0[1560] | layer_0[1015]); 
    assign out[421] = ~layer_0[85]; 
    assign out[422] = layer_0[2377] ^ layer_0[1031]; 
    assign out[423] = ~layer_0[1563]; 
    assign out[424] = layer_0[241] | layer_0[808]; 
    assign out[425] = ~(layer_0[683] ^ layer_0[1017]); 
    assign out[426] = layer_0[838] ^ layer_0[1230]; 
    assign out[427] = ~(layer_0[2528] | layer_0[28]); 
    assign out[428] = layer_0[2507] | layer_0[15]; 
    assign out[429] = ~(layer_0[1866] ^ layer_0[1340]); 
    assign out[430] = layer_0[283] & ~layer_0[2450]; 
    assign out[431] = layer_0[1975] & ~layer_0[883]; 
    assign out[432] = ~(layer_0[1370] ^ layer_0[1778]); 
    assign out[433] = layer_0[185] & ~layer_0[2184]; 
    assign out[434] = layer_0[251] & ~layer_0[1775]; 
    assign out[435] = layer_0[1868] & ~layer_0[1797]; 
    assign out[436] = layer_0[1861]; 
    assign out[437] = ~(layer_0[1887] ^ layer_0[92]); 
    assign out[438] = ~layer_0[1577]; 
    assign out[439] = layer_0[2486] & layer_0[931]; 
    assign out[440] = ~layer_0[2287]; 
    assign out[441] = layer_0[1699] ^ layer_0[102]; 
    assign out[442] = ~layer_0[2491]; 
    assign out[443] = layer_0[1604] | layer_0[0]; 
    assign out[444] = ~(layer_0[1914] | layer_0[2120]); 
    assign out[445] = layer_0[1791]; 
    assign out[446] = ~(layer_0[1809] | layer_0[1778]); 
    assign out[447] = ~(layer_0[219] | layer_0[809]); 
    assign out[448] = ~(layer_0[8] ^ layer_0[2244]); 
    assign out[449] = layer_0[1985]; 
    assign out[450] = ~(layer_0[766] & layer_0[1958]); 
    assign out[451] = layer_0[294]; 
    assign out[452] = ~(layer_0[1913] | layer_0[696]); 
    assign out[453] = layer_0[2520] ^ layer_0[2352]; 
    assign out[454] = layer_0[1641] & ~layer_0[1900]; 
    assign out[455] = ~(layer_0[176] | layer_0[1751]); 
    assign out[456] = layer_0[765] ^ layer_0[567]; 
    assign out[457] = layer_0[1022] & ~layer_0[650]; 
    assign out[458] = ~layer_0[1560]; 
    assign out[459] = layer_0[1654] & layer_0[1791]; 
    assign out[460] = layer_0[931] & ~layer_0[1251]; 
    assign out[461] = layer_0[2282] & layer_0[601]; 
    assign out[462] = ~(layer_0[1966] ^ layer_0[2406]); 
    assign out[463] = ~(layer_0[665] | layer_0[2316]); 
    assign out[464] = ~layer_0[1111]; 
    assign out[465] = layer_0[2286] & ~layer_0[1971]; 
    assign out[466] = ~(layer_0[2069] | layer_0[2288]); 
    assign out[467] = ~(layer_0[1351] ^ layer_0[111]); 
    assign out[468] = layer_0[1196] ^ layer_0[1509]; 
    assign out[469] = layer_0[1044] & layer_0[1856]; 
    assign out[470] = layer_0[2267] & ~layer_0[651]; 
    assign out[471] = layer_0[1389] & ~layer_0[440]; 
    assign out[472] = ~(layer_0[1325] ^ layer_0[1470]); 
    assign out[473] = layer_0[31] ^ layer_0[486]; 
    assign out[474] = ~(layer_0[482] ^ layer_0[1592]); 
    assign out[475] = layer_0[1596]; 
    assign out[476] = layer_0[202]; 
    assign out[477] = layer_0[49] & ~layer_0[1860]; 
    assign out[478] = layer_0[1247]; 
    assign out[479] = layer_0[1109] ^ layer_0[1735]; 
    assign out[480] = layer_0[352] & ~layer_0[686]; 
    assign out[481] = ~(layer_0[2169] ^ layer_0[1109]); 
    assign out[482] = layer_0[612]; 
    assign out[483] = ~(layer_0[1703] ^ layer_0[383]); 
    assign out[484] = ~(layer_0[543] ^ layer_0[2202]); 
    assign out[485] = layer_0[1821] ^ layer_0[2152]; 
    assign out[486] = layer_0[870]; 
    assign out[487] = layer_0[1604] ^ layer_0[1097]; 
    assign out[488] = ~(layer_0[492] ^ layer_0[62]); 
    assign out[489] = layer_0[1963] & layer_0[846]; 
    assign out[490] = layer_0[1256] ^ layer_0[349]; 
    assign out[491] = layer_0[320] & ~layer_0[1229]; 
    assign out[492] = layer_0[349] & ~layer_0[1705]; 
    assign out[493] = ~(layer_0[2025] ^ layer_0[387]); 
    assign out[494] = ~(layer_0[1463] ^ layer_0[2504]); 
    assign out[495] = ~(layer_0[1660] ^ layer_0[526]); 
    assign out[496] = ~layer_0[1556]; 
    assign out[497] = ~layer_0[1670] | (layer_0[1552] & layer_0[1670]); 
    assign out[498] = layer_0[487] & ~layer_0[63]; 
    assign out[499] = layer_0[1580] & ~layer_0[1209]; 
    assign out[500] = ~layer_0[1873]; 
    assign out[501] = layer_0[2213]; 
    assign out[502] = ~(layer_0[1767] ^ layer_0[1019]); 
    assign out[503] = layer_0[1794] & layer_0[606]; 
    assign out[504] = layer_0[312] ^ layer_0[888]; 
    assign out[505] = layer_0[113] ^ layer_0[2295]; 
    assign out[506] = ~layer_0[565]; 
    assign out[507] = ~layer_0[2531]; 
    assign out[508] = layer_0[1652] & ~layer_0[176]; 
    assign out[509] = ~(layer_0[1774] ^ layer_0[1693]); 
    assign out[510] = layer_0[470]; 
    assign out[511] = layer_0[2026] | layer_0[1070]; 
    assign out[512] = ~(layer_0[147] ^ layer_0[906]); 
    assign out[513] = ~(layer_0[2080] & layer_0[257]); 
    assign out[514] = ~(layer_0[1319] ^ layer_0[1424]); 
    assign out[515] = ~(layer_0[300] | layer_0[1578]); 
    assign out[516] = ~(layer_0[1534] ^ layer_0[1141]); 
    assign out[517] = ~layer_0[1719]; 
    assign out[518] = layer_0[425]; 
    assign out[519] = ~(layer_0[2030] ^ layer_0[702]); 
    assign out[520] = layer_0[1881] & ~layer_0[797]; 
    assign out[521] = ~layer_0[928] | (layer_0[928] & layer_0[2159]); 
    assign out[522] = layer_0[2223] ^ layer_0[1413]; 
    assign out[523] = layer_0[1381] ^ layer_0[612]; 
    assign out[524] = ~(layer_0[1499] ^ layer_0[841]); 
    assign out[525] = ~layer_0[1801]; 
    assign out[526] = layer_0[1884] & ~layer_0[1898]; 
    assign out[527] = layer_0[811]; 
    assign out[528] = ~layer_0[101]; 
    assign out[529] = layer_0[1193] & ~layer_0[580]; 
    assign out[530] = ~(layer_0[2226] ^ layer_0[2333]); 
    assign out[531] = ~(layer_0[980] & layer_0[1217]); 
    assign out[532] = ~(layer_0[1852] ^ layer_0[2251]); 
    assign out[533] = layer_0[1868] & ~layer_0[2024]; 
    assign out[534] = ~layer_0[48]; 
    assign out[535] = layer_0[1110]; 
    assign out[536] = layer_0[1906] & layer_0[1816]; 
    assign out[537] = layer_0[1990] ^ layer_0[2403]; 
    assign out[538] = layer_0[1691] | layer_0[1295]; 
    assign out[539] = layer_0[771]; 
    assign out[540] = ~(layer_0[1602] ^ layer_0[1892]); 
    assign out[541] = ~layer_0[2349]; 
    assign out[542] = ~layer_0[1750] | (layer_0[2510] & layer_0[1750]); 
    assign out[543] = layer_0[674]; 
    assign out[544] = ~layer_0[1808]; 
    assign out[545] = ~(layer_0[1887] ^ layer_0[1143]); 
    assign out[546] = layer_0[425]; 
    assign out[547] = ~layer_0[2360]; 
    assign out[548] = ~layer_0[76] | (layer_0[1954] & layer_0[76]); 
    assign out[549] = layer_0[1757] ^ layer_0[450]; 
    assign out[550] = layer_0[1746] ^ layer_0[2439]; 
    assign out[551] = ~layer_0[715]; 
    assign out[552] = layer_0[1963] ^ layer_0[1567]; 
    assign out[553] = layer_0[408] ^ layer_0[2313]; 
    assign out[554] = layer_0[754] & ~layer_0[1551]; 
    assign out[555] = ~(layer_0[1472] ^ layer_0[1262]); 
    assign out[556] = layer_0[445]; 
    assign out[557] = layer_0[1868]; 
    assign out[558] = layer_0[522] & ~layer_0[810]; 
    assign out[559] = layer_0[470] & ~layer_0[95]; 
    assign out[560] = ~layer_0[333]; 
    assign out[561] = layer_0[1427] ^ layer_0[1650]; 
    assign out[562] = ~(layer_0[2025] | layer_0[411]); 
    assign out[563] = layer_0[2056] & ~layer_0[1902]; 
    assign out[564] = layer_0[2068] ^ layer_0[954]; 
    assign out[565] = ~(layer_0[1670] ^ layer_0[2157]); 
    assign out[566] = layer_0[701] | layer_0[1923]; 
    assign out[567] = ~(layer_0[505] ^ layer_0[2042]); 
    assign out[568] = ~(layer_0[1124] & layer_0[1456]); 
    assign out[569] = ~(layer_0[2463] & layer_0[2421]); 
    assign out[570] = layer_0[374] ^ layer_0[1376]; 
    assign out[571] = ~layer_0[882]; 
    assign out[572] = layer_0[555] | layer_0[1616]; 
    assign out[573] = ~(layer_0[991] ^ layer_0[154]); 
    assign out[574] = layer_0[2038] & ~layer_0[2084]; 
    assign out[575] = ~layer_0[605] | (layer_0[1450] & layer_0[605]); 
    assign out[576] = layer_0[441] | layer_0[88]; 
    assign out[577] = layer_0[881]; 
    assign out[578] = layer_0[1816]; 
    assign out[579] = ~layer_0[882]; 
    assign out[580] = ~(layer_0[2395] ^ layer_0[570]); 
    assign out[581] = layer_0[2304] ^ layer_0[57]; 
    assign out[582] = layer_0[966] & ~layer_0[101]; 
    assign out[583] = ~layer_0[1270]; 
    assign out[584] = ~layer_0[2001] | (layer_0[2001] & layer_0[401]); 
    assign out[585] = layer_0[336]; 
    assign out[586] = ~(layer_0[2333] ^ layer_0[997]); 
    assign out[587] = ~layer_0[1200]; 
    assign out[588] = layer_0[1379] ^ layer_0[294]; 
    assign out[589] = layer_0[2282] & ~layer_0[2087]; 
    assign out[590] = ~(layer_0[2408] ^ layer_0[1784]); 
    assign out[591] = layer_0[558]; 
    assign out[592] = ~(layer_0[1735] & layer_0[1411]); 
    assign out[593] = layer_0[754] ^ layer_0[605]; 
    assign out[594] = layer_0[555]; 
    assign out[595] = ~(layer_0[2301] | layer_0[373]); 
    assign out[596] = ~(layer_0[750] ^ layer_0[1960]); 
    assign out[597] = layer_0[113] ^ layer_0[1830]; 
    assign out[598] = layer_0[2510] | layer_0[856]; 
    assign out[599] = ~(layer_0[1017] | layer_0[2207]); 
    assign out[600] = layer_0[680] & ~layer_0[67]; 
    assign out[601] = ~(layer_0[1229] ^ layer_0[160]); 
    assign out[602] = layer_0[2230]; 
    assign out[603] = ~(layer_0[2393] | layer_0[301]); 
    assign out[604] = ~layer_0[1818]; 
    assign out[605] = ~(layer_0[329] ^ layer_0[552]); 
    assign out[606] = ~layer_0[357] | (layer_0[357] & layer_0[2026]); 
    assign out[607] = layer_0[202]; 
    assign out[608] = layer_0[1194] ^ layer_0[1588]; 
    assign out[609] = ~layer_0[960]; 
    assign out[610] = ~(layer_0[520] ^ layer_0[739]); 
    assign out[611] = layer_0[327]; 
    assign out[612] = layer_0[160]; 
    assign out[613] = ~layer_0[980] | (layer_0[980] & layer_0[712]); 
    assign out[614] = layer_0[463] ^ layer_0[2061]; 
    assign out[615] = layer_0[2454] & layer_0[1075]; 
    assign out[616] = layer_0[2056]; 
    assign out[617] = layer_0[1118] & ~layer_0[1366]; 
    assign out[618] = ~(layer_0[764] | layer_0[2536]); 
    assign out[619] = ~layer_0[1306] | (layer_0[1306] & layer_0[919]); 
    assign out[620] = layer_0[2221]; 
    assign out[621] = ~(layer_0[1750] & layer_0[1157]); 
    assign out[622] = layer_0[1941]; 
    assign out[623] = layer_0[1840] ^ layer_0[1580]; 
    assign out[624] = ~layer_0[84] | (layer_0[84] & layer_0[1700]); 
    assign out[625] = layer_0[555] & ~layer_0[606]; 
    assign out[626] = ~(layer_0[2246] ^ layer_0[1867]); 
    assign out[627] = ~(layer_0[1489] | layer_0[2340]); 
    assign out[628] = ~layer_0[2181]; 
    assign out[629] = ~layer_0[1178]; 
    assign out[630] = ~layer_0[411] | (layer_0[145] & layer_0[411]); 
    assign out[631] = ~(layer_0[360] ^ layer_0[1241]); 
    assign out[632] = ~layer_0[1139]; 
    assign out[633] = ~(layer_0[878] ^ layer_0[382]); 
    assign out[634] = layer_0[1900]; 
    assign out[635] = layer_0[1954] & layer_0[1150]; 
    assign out[636] = layer_0[1942] ^ layer_0[1704]; 
    assign out[637] = ~(layer_0[2251] | layer_0[2156]); 
    assign out[638] = ~layer_0[1853]; 
    assign out[639] = layer_0[1450] & layer_0[1746]; 
    assign out[640] = ~(layer_0[531] ^ layer_0[1625]); 
    assign out[641] = layer_0[1209] ^ layer_0[514]; 
    assign out[642] = layer_0[2038]; 
    assign out[643] = ~(layer_0[2485] ^ layer_0[1459]); 
    assign out[644] = layer_0[1690] & ~layer_0[863]; 
    assign out[645] = ~layer_0[1995]; 
    assign out[646] = ~(layer_0[1872] | layer_0[715]); 
    assign out[647] = ~(layer_0[151] ^ layer_0[1712]); 
    assign out[648] = layer_0[131] ^ layer_0[1367]; 
    assign out[649] = layer_0[1770] ^ layer_0[1245]; 
    assign out[650] = layer_0[5] & ~layer_0[2351]; 
    assign out[651] = layer_0[272] ^ layer_0[323]; 
    assign out[652] = layer_0[1557] ^ layer_0[1422]; 
    assign out[653] = ~layer_0[2049] | (layer_0[558] & layer_0[2049]); 
    assign out[654] = layer_0[2077] ^ layer_0[1250]; 
    assign out[655] = ~(layer_0[1265] ^ layer_0[1157]); 
    assign out[656] = ~(layer_0[2492] & layer_0[1548]); 
    assign out[657] = ~(layer_0[716] ^ layer_0[123]); 
    assign out[658] = layer_0[2199]; 
    assign out[659] = layer_0[400] ^ layer_0[2200]; 
    assign out[660] = ~layer_0[101]; 
    assign out[661] = ~layer_0[2162]; 
    assign out[662] = layer_0[99]; 
    assign out[663] = layer_0[2266] ^ layer_0[555]; 
    assign out[664] = ~(layer_0[486] ^ layer_0[2436]); 
    assign out[665] = layer_0[733]; 
    assign out[666] = ~(layer_0[853] ^ layer_0[1244]); 
    assign out[667] = ~layer_0[448]; 
    assign out[668] = ~layer_0[1898] | (layer_0[1473] & layer_0[1898]); 
    assign out[669] = ~(layer_0[1439] | layer_0[1416]); 
    assign out[670] = layer_0[919] ^ layer_0[517]; 
    assign out[671] = ~(layer_0[992] | layer_0[1054]); 
    assign out[672] = layer_0[1091] | layer_0[799]; 
    assign out[673] = layer_0[572]; 
    assign out[674] = layer_0[1813] | layer_0[174]; 
    assign out[675] = layer_0[1977] ^ layer_0[1699]; 
    assign out[676] = layer_0[672] ^ layer_0[206]; 
    assign out[677] = ~layer_0[1995]; 
    assign out[678] = layer_0[476] ^ layer_0[775]; 
    assign out[679] = ~layer_0[694]; 
    assign out[680] = layer_0[123] & ~layer_0[1924]; 
    assign out[681] = ~(layer_0[2053] & layer_0[127]); 
    assign out[682] = layer_0[1584] & ~layer_0[210]; 
    assign out[683] = ~(layer_0[2046] | layer_0[1173]); 
    assign out[684] = ~(layer_0[1528] ^ layer_0[989]); 
    assign out[685] = ~(layer_0[1291] | layer_0[380]); 
    assign out[686] = layer_0[1523] ^ layer_0[2072]; 
    assign out[687] = ~layer_0[2083] | (layer_0[1813] & layer_0[2083]); 
    assign out[688] = ~layer_0[696] | (layer_0[696] & layer_0[627]); 
    assign out[689] = ~(layer_0[980] ^ layer_0[966]); 
    assign out[690] = layer_0[1404]; 
    assign out[691] = ~layer_0[378] | (layer_0[378] & layer_0[2542]); 
    assign out[692] = ~layer_0[1788] | (layer_0[1788] & layer_0[1261]); 
    assign out[693] = layer_0[2077]; 
    assign out[694] = ~layer_0[67]; 
    assign out[695] = ~(layer_0[1518] | layer_0[1397]); 
    assign out[696] = layer_0[1633]; 
    assign out[697] = ~(layer_0[2221] ^ layer_0[1236]); 
    assign out[698] = layer_0[2178] ^ layer_0[929]; 
    assign out[699] = layer_0[353]; 
    assign out[700] = ~layer_0[1181]; 
    assign out[701] = layer_0[100] | layer_0[201]; 
    assign out[702] = layer_0[2348] | layer_0[1827]; 
    assign out[703] = layer_0[1260] & ~layer_0[1522]; 
    assign out[704] = ~layer_0[1180]; 
    assign out[705] = ~layer_0[1621] | (layer_0[1477] & layer_0[1621]); 
    assign out[706] = layer_0[1828] ^ layer_0[213]; 
    assign out[707] = layer_0[538] & layer_0[1167]; 
    assign out[708] = ~layer_0[1274]; 
    assign out[709] = layer_0[1262]; 
    assign out[710] = layer_0[1428]; 
    assign out[711] = ~layer_0[1578] | (layer_0[1862] & layer_0[1578]); 
    assign out[712] = ~(layer_0[2024] ^ layer_0[1920]); 
    assign out[713] = layer_0[160]; 
    assign out[714] = layer_0[412] & ~layer_0[609]; 
    assign out[715] = ~layer_0[210]; 
    assign out[716] = ~(layer_0[1451] ^ layer_0[1536]); 
    assign out[717] = layer_0[2310] & layer_0[61]; 
    assign out[718] = ~(layer_0[1356] | layer_0[2407]); 
    assign out[719] = ~(layer_0[395] ^ layer_0[2006]); 
    assign out[720] = ~layer_0[943]; 
    assign out[721] = layer_0[467] ^ layer_0[1877]; 
    assign out[722] = ~layer_0[140]; 
    assign out[723] = layer_0[1906]; 
    assign out[724] = layer_0[123] & layer_0[811]; 
    assign out[725] = layer_0[485] ^ layer_0[1162]; 
    assign out[726] = layer_0[2089] & ~layer_0[1403]; 
    assign out[727] = ~layer_0[67]; 
    assign out[728] = ~layer_0[2162]; 
    assign out[729] = layer_0[99] & ~layer_0[2254]; 
    assign out[730] = ~(layer_0[380] ^ layer_0[1486]); 
    assign out[731] = layer_0[1848]; 
    assign out[732] = ~(layer_0[267] ^ layer_0[1027]); 
    assign out[733] = ~(layer_0[2219] ^ layer_0[1686]); 
    assign out[734] = ~(layer_0[2207] | layer_0[300]); 
    assign out[735] = ~layer_0[1333] | (layer_0[1388] & layer_0[1333]); 
    assign out[736] = ~layer_0[847]; 
    assign out[737] = layer_0[1401] ^ layer_0[2101]; 
    assign out[738] = layer_0[1472]; 
    assign out[739] = layer_0[2531]; 
    assign out[740] = ~layer_0[155] | (layer_0[155] & layer_0[458]); 
    assign out[741] = layer_0[286]; 
    assign out[742] = layer_0[332] | layer_0[2329]; 
    assign out[743] = ~(layer_0[2405] ^ layer_0[427]); 
    assign out[744] = layer_0[885] ^ layer_0[1110]; 
    assign out[745] = layer_0[184] ^ layer_0[650]; 
    assign out[746] = ~layer_0[1374] | (layer_0[1374] & layer_0[1076]); 
    assign out[747] = ~(layer_0[2257] | layer_0[2249]); 
    assign out[748] = layer_0[1897] ^ layer_0[876]; 
    assign out[749] = ~layer_0[585] | (layer_0[585] & layer_0[2242]); 
    assign out[750] = ~layer_0[1836]; 
    assign out[751] = layer_0[1230] ^ layer_0[1143]; 
    assign out[752] = layer_0[881]; 
    assign out[753] = layer_0[2252] & ~layer_0[2372]; 
    assign out[754] = layer_0[174]; 
    assign out[755] = ~(layer_0[318] | layer_0[2181]); 
    assign out[756] = ~layer_0[95]; 
    assign out[757] = layer_0[741]; 
    assign out[758] = layer_0[2242] & ~layer_0[2437]; 
    assign out[759] = ~(layer_0[1727] ^ layer_0[729]); 
    assign out[760] = layer_0[1522] ^ layer_0[1743]; 
    assign out[761] = ~layer_0[63] | (layer_0[63] & layer_0[632]); 
    assign out[762] = ~layer_0[1157]; 
    assign out[763] = ~(layer_0[2099] ^ layer_0[1297]); 
    assign out[764] = layer_0[313]; 
    assign out[765] = layer_0[2039]; 
    assign out[766] = ~layer_0[689]; 
    assign out[767] = ~layer_0[1141]; 
    assign out[768] = layer_0[1346] ^ layer_0[852]; 
    assign out[769] = layer_0[652] ^ layer_0[375]; 
    assign out[770] = ~(layer_0[805] | layer_0[2517]); 
    assign out[771] = layer_0[1057] & layer_0[821]; 
    assign out[772] = layer_0[1020] ^ layer_0[1699]; 
    assign out[773] = layer_0[378] & layer_0[2458]; 
    assign out[774] = layer_0[1143] ^ layer_0[1043]; 
    assign out[775] = layer_0[2324] & ~layer_0[1069]; 
    assign out[776] = ~(layer_0[1593] ^ layer_0[2533]); 
    assign out[777] = layer_0[1908] & ~layer_0[1297]; 
    assign out[778] = ~(layer_0[2212] ^ layer_0[173]); 
    assign out[779] = layer_0[663]; 
    assign out[780] = ~(layer_0[1516] | layer_0[1003]); 
    assign out[781] = layer_0[2149]; 
    assign out[782] = layer_0[1886] | layer_0[2227]; 
    assign out[783] = layer_0[1292] ^ layer_0[1439]; 
    assign out[784] = layer_0[1399] & ~layer_0[1107]; 
    assign out[785] = ~layer_0[2354] | (layer_0[2354] & layer_0[242]); 
    assign out[786] = ~(layer_0[2376] ^ layer_0[1798]); 
    assign out[787] = layer_0[1073] ^ layer_0[834]; 
    assign out[788] = layer_0[1762] & layer_0[557]; 
    assign out[789] = layer_0[485] ^ layer_0[2525]; 
    assign out[790] = ~(layer_0[355] ^ layer_0[1030]); 
    assign out[791] = layer_0[96] & ~layer_0[2055]; 
    assign out[792] = ~layer_0[2226]; 
    assign out[793] = ~layer_0[599]; 
    assign out[794] = ~layer_0[2368]; 
    assign out[795] = layer_0[393]; 
    assign out[796] = layer_0[393] ^ layer_0[287]; 
    assign out[797] = ~layer_0[1352]; 
    assign out[798] = ~layer_0[1503] | (layer_0[128] & layer_0[1503]); 
    assign out[799] = ~(layer_0[1004] ^ layer_0[1654]); 
    assign out[800] = layer_0[2102] & layer_0[1022]; 
    assign out[801] = ~layer_0[620]; 
    assign out[802] = ~(layer_0[2518] | layer_0[1444]); 
    assign out[803] = ~(layer_0[994] ^ layer_0[267]); 
    assign out[804] = ~(layer_0[221] ^ layer_0[2507]); 
    assign out[805] = ~(layer_0[1619] ^ layer_0[1028]); 
    assign out[806] = ~layer_0[1184]; 
    assign out[807] = layer_0[1484]; 
    assign out[808] = ~layer_0[161]; 
    assign out[809] = layer_0[1393] ^ layer_0[1686]; 
    assign out[810] = ~layer_0[2196] | (layer_0[2196] & layer_0[912]); 
    assign out[811] = layer_0[2523] ^ layer_0[144]; 
    assign out[812] = ~layer_0[1025]; 
    assign out[813] = ~layer_0[753]; 
    assign out[814] = layer_0[2053]; 
    assign out[815] = layer_0[2379] & layer_0[1137]; 
    assign out[816] = layer_0[2404] & layer_0[2042]; 
    assign out[817] = ~layer_0[1857] | (layer_0[1857] & layer_0[638]); 
    assign out[818] = layer_0[1495] & ~layer_0[2253]; 
    assign out[819] = ~(layer_0[1090] ^ layer_0[1819]); 
    assign out[820] = layer_0[1799] ^ layer_0[8]; 
    assign out[821] = layer_0[1828] & ~layer_0[1357]; 
    assign out[822] = layer_0[2142]; 
    assign out[823] = layer_0[479] & ~layer_0[1851]; 
    assign out[824] = ~(layer_0[2300] ^ layer_0[751]); 
    assign out[825] = ~layer_0[2340]; 
    assign out[826] = layer_0[173]; 
    assign out[827] = ~layer_0[1256] | (layer_0[1256] & layer_0[530]); 
    assign out[828] = ~(layer_0[914] ^ layer_0[2138]); 
    assign out[829] = ~layer_0[495]; 
    assign out[830] = layer_0[1262] & ~layer_0[1129]; 
    assign out[831] = layer_0[1908]; 
    assign out[832] = ~(layer_0[2552] ^ layer_0[165]); 
    assign out[833] = layer_0[288] & layer_0[348]; 
    assign out[834] = ~layer_0[1357]; 
    assign out[835] = ~layer_0[995]; 
    assign out[836] = ~(layer_0[1690] ^ layer_0[2258]); 
    assign out[837] = ~layer_0[62] | (layer_0[1855] & layer_0[62]); 
    assign out[838] = layer_0[1155] & ~layer_0[1996]; 
    assign out[839] = ~layer_0[1823] | (layer_0[1823] & layer_0[2396]); 
    assign out[840] = layer_0[496]; 
    assign out[841] = ~layer_0[310] | (layer_0[310] & layer_0[1852]); 
    assign out[842] = layer_0[2142]; 
    assign out[843] = layer_0[417] & layer_0[1721]; 
    assign out[844] = layer_0[1367] ^ layer_0[413]; 
    assign out[845] = ~layer_0[1919]; 
    assign out[846] = layer_0[266]; 
    assign out[847] = ~layer_0[1283]; 
    assign out[848] = ~layer_0[711] | (layer_0[744] & layer_0[711]); 
    assign out[849] = layer_0[1077] & ~layer_0[1593]; 
    assign out[850] = layer_0[1081] | layer_0[198]; 
    assign out[851] = layer_0[1448]; 
    assign out[852] = ~(layer_0[208] ^ layer_0[515]); 
    assign out[853] = layer_0[117] ^ layer_0[1677]; 
    assign out[854] = ~(layer_0[392] & layer_0[411]); 
    assign out[855] = ~layer_0[676]; 
    assign out[856] = layer_0[203] ^ layer_0[1251]; 
    assign out[857] = layer_0[2268] & layer_0[2022]; 
    assign out[858] = ~layer_0[2050] | (layer_0[2050] & layer_0[903]); 
    assign out[859] = layer_0[879] | layer_0[2176]; 
    assign out[860] = layer_0[2301]; 
    assign out[861] = layer_0[2225] & ~layer_0[2067]; 
    assign out[862] = layer_0[2487] & ~layer_0[641]; 
    assign out[863] = ~layer_0[1547]; 
    assign out[864] = ~(layer_0[262] ^ layer_0[2303]); 
    assign out[865] = layer_0[662] & ~layer_0[1587]; 
    assign out[866] = layer_0[977] ^ layer_0[1994]; 
    assign out[867] = layer_0[524]; 
    assign out[868] = ~layer_0[1197]; 
    assign out[869] = ~(layer_0[412] | layer_0[1735]); 
    assign out[870] = layer_0[815]; 
    assign out[871] = ~layer_0[106]; 
    assign out[872] = layer_0[706] & ~layer_0[484]; 
    assign out[873] = ~(layer_0[1107] & layer_0[2392]); 
    assign out[874] = ~layer_0[1023] | (layer_0[1023] & layer_0[479]); 
    assign out[875] = ~(layer_0[499] | layer_0[586]); 
    assign out[876] = layer_0[181]; 
    assign out[877] = ~(layer_0[133] ^ layer_0[1859]); 
    assign out[878] = layer_0[9] & layer_0[1262]; 
    assign out[879] = layer_0[370]; 
    assign out[880] = ~(layer_0[2423] ^ layer_0[2302]); 
    assign out[881] = ~(layer_0[1769] ^ layer_0[2009]); 
    assign out[882] = layer_0[553]; 
    assign out[883] = ~(layer_0[1348] & layer_0[1739]); 
    assign out[884] = ~layer_0[705]; 
    assign out[885] = layer_0[201] & layer_0[1838]; 
    assign out[886] = layer_0[395] & ~layer_0[1716]; 
    assign out[887] = ~(layer_0[899] ^ layer_0[1459]); 
    assign out[888] = layer_0[2427] & layer_0[269]; 
    assign out[889] = ~(layer_0[2112] ^ layer_0[1542]); 
    assign out[890] = ~layer_0[2158]; 
    assign out[891] = ~layer_0[1655]; 
    assign out[892] = layer_0[2298]; 
    assign out[893] = ~layer_0[1353] | (layer_0[1353] & layer_0[395]); 
    assign out[894] = ~layer_0[1293]; 
    assign out[895] = layer_0[224] ^ layer_0[833]; 
    assign out[896] = ~(layer_0[1050] ^ layer_0[310]); 
    assign out[897] = layer_0[1260]; 
    assign out[898] = ~(layer_0[1263] ^ layer_0[1574]); 
    assign out[899] = ~layer_0[244]; 
    assign out[900] = ~(layer_0[920] | layer_0[36]); 
    assign out[901] = ~layer_0[724]; 
    assign out[902] = layer_0[1042] & ~layer_0[1283]; 
    assign out[903] = layer_0[242] | layer_0[1132]; 
    assign out[904] = layer_0[2379] & ~layer_0[0]; 
    assign out[905] = layer_0[888]; 
    assign out[906] = layer_0[2388] & layer_0[911]; 
    assign out[907] = layer_0[416] ^ layer_0[395]; 
    assign out[908] = ~(layer_0[655] | layer_0[1537]); 
    assign out[909] = layer_0[1828] & layer_0[2136]; 
    assign out[910] = ~layer_0[1394]; 
    assign out[911] = ~layer_0[1537] | (layer_0[1342] & layer_0[1537]); 
    assign out[912] = ~(layer_0[920] ^ layer_0[308]); 
    assign out[913] = ~layer_0[664]; 
    assign out[914] = layer_0[948]; 
    assign out[915] = layer_0[227]; 
    assign out[916] = layer_0[1354] & ~layer_0[1534]; 
    assign out[917] = ~layer_0[1214]; 
    assign out[918] = layer_0[1623] ^ layer_0[1891]; 
    assign out[919] = layer_0[1046] ^ layer_0[1630]; 
    assign out[920] = layer_0[404] ^ layer_0[394]; 
    assign out[921] = ~(layer_0[1629] | layer_0[2076]); 
    assign out[922] = layer_0[2482] & ~layer_0[1629]; 
    assign out[923] = layer_0[2051]; 
    assign out[924] = layer_0[2149] & ~layer_0[428]; 
    assign out[925] = layer_0[1697] ^ layer_0[1426]; 
    assign out[926] = layer_0[2219]; 
    assign out[927] = ~layer_0[1033]; 
    assign out[928] = ~(layer_0[1367] ^ layer_0[1924]); 
    assign out[929] = layer_0[1576]; 
    assign out[930] = layer_0[2302]; 
    assign out[931] = layer_0[564] ^ layer_0[2267]; 
    assign out[932] = ~(layer_0[1048] ^ layer_0[2262]); 
    assign out[933] = ~(layer_0[383] ^ layer_0[284]); 
    assign out[934] = ~(layer_0[1346] | layer_0[1804]); 
    assign out[935] = layer_0[2009] ^ layer_0[931]; 
    assign out[936] = ~layer_0[1104]; 
    assign out[937] = ~layer_0[1914]; 
    assign out[938] = layer_0[826] ^ layer_0[1407]; 
    assign out[939] = ~layer_0[2167] | (layer_0[2167] & layer_0[982]); 
    assign out[940] = layer_0[989] ^ layer_0[1576]; 
    assign out[941] = ~layer_0[594]; 
    assign out[942] = ~(layer_0[1661] ^ layer_0[1782]); 
    assign out[943] = layer_0[2053]; 
    assign out[944] = layer_0[1354] & layer_0[1923]; 
    assign out[945] = layer_0[646]; 
    assign out[946] = ~layer_0[532]; 
    assign out[947] = layer_0[1516] ^ layer_0[1494]; 
    assign out[948] = ~layer_0[901]; 
    assign out[949] = ~(layer_0[1317] | layer_0[1820]); 
    assign out[950] = ~layer_0[384] | (layer_0[384] & layer_0[194]); 
    assign out[951] = layer_0[539] ^ layer_0[2405]; 
    assign out[952] = layer_0[1675]; 
    assign out[953] = ~(layer_0[511] ^ layer_0[1976]); 
    assign out[954] = layer_0[2168] ^ layer_0[468]; 
    assign out[955] = layer_0[577] & ~layer_0[1877]; 
    assign out[956] = layer_0[1048] ^ layer_0[1327]; 
    assign out[957] = layer_0[445] & ~layer_0[591]; 
    assign out[958] = layer_0[765] & ~layer_0[2328]; 
    assign out[959] = layer_0[488]; 
    assign out[960] = ~layer_0[664]; 
    assign out[961] = ~layer_0[2400]; 
    assign out[962] = layer_0[1483] ^ layer_0[937]; 
    assign out[963] = ~layer_0[274]; 
    assign out[964] = layer_0[1511] ^ layer_0[1745]; 
    assign out[965] = layer_0[1541] & ~layer_0[280]; 
    assign out[966] = layer_0[779] ^ layer_0[1918]; 
    assign out[967] = layer_0[2537] ^ layer_0[2493]; 
    assign out[968] = ~(layer_0[699] ^ layer_0[271]); 
    assign out[969] = layer_0[305]; 
    assign out[970] = ~(layer_0[627] | layer_0[1069]); 
    assign out[971] = layer_0[194]; 
    assign out[972] = ~layer_0[2384]; 
    assign out[973] = layer_0[1949] ^ layer_0[2022]; 
    assign out[974] = layer_0[964] & ~layer_0[1692]; 
    assign out[975] = layer_0[559] & ~layer_0[689]; 
    assign out[976] = ~layer_0[2110]; 
    assign out[977] = layer_0[377] & ~layer_0[1069]; 
    assign out[978] = layer_0[2388]; 
    assign out[979] = layer_0[2218] & ~layer_0[1357]; 
    assign out[980] = ~(layer_0[2061] ^ layer_0[1316]); 
    assign out[981] = layer_0[309] | layer_0[1509]; 
    assign out[982] = ~layer_0[134]; 
    assign out[983] = ~(layer_0[549] ^ layer_0[544]); 
    assign out[984] = layer_0[1243] ^ layer_0[220]; 
    assign out[985] = ~layer_0[932]; 
    assign out[986] = layer_0[761] ^ layer_0[1318]; 
    assign out[987] = layer_0[210] ^ layer_0[888]; 
    assign out[988] = layer_0[1226] & layer_0[22]; 
    assign out[989] = ~layer_0[1450]; 
    assign out[990] = ~layer_0[1558]; 
    assign out[991] = ~layer_0[901] | (layer_0[901] & layer_0[206]); 
    assign out[992] = layer_0[1203] ^ layer_0[954]; 
    assign out[993] = layer_0[1764]; 
    assign out[994] = ~(layer_0[968] ^ layer_0[1112]); 
    assign out[995] = layer_0[1006] & layer_0[2260]; 
    assign out[996] = ~(layer_0[1930] | layer_0[2078]); 
    assign out[997] = layer_0[1613] & layer_0[127]; 
    assign out[998] = layer_0[209]; 
    assign out[999] = ~layer_0[121]; 
    assign out[1000] = ~(layer_0[1802] ^ layer_0[1371]); 
    assign out[1001] = layer_0[1490] & ~layer_0[2414]; 
    assign out[1002] = ~layer_0[1379] | (layer_0[1056] & layer_0[1379]); 
    assign out[1003] = layer_0[479]; 
    assign out[1004] = ~(layer_0[2303] | layer_0[2173]); 
    assign out[1005] = ~layer_0[2128]; 
    assign out[1006] = layer_0[798] & ~layer_0[2201]; 
    assign out[1007] = ~layer_0[907] | (layer_0[907] & layer_0[2396]); 
    assign out[1008] = ~layer_0[121]; 
    assign out[1009] = ~(layer_0[1498] ^ layer_0[184]); 
    assign out[1010] = ~(layer_0[731] | layer_0[2400]); 
    assign out[1011] = ~layer_0[441] | (layer_0[1682] & layer_0[441]); 
    assign out[1012] = layer_0[1229] ^ layer_0[2267]; 
    assign out[1013] = layer_0[31] ^ layer_0[818]; 
    assign out[1014] = ~(layer_0[11] ^ layer_0[1548]); 
    assign out[1015] = layer_0[652] ^ layer_0[1926]; 
    assign out[1016] = layer_0[1937] ^ layer_0[1529]; 
    assign out[1017] = layer_0[52]; 
    assign out[1018] = ~(layer_0[2228] | layer_0[2400]); 
    assign out[1019] = ~(layer_0[1795] ^ layer_0[350]); 
    assign out[1020] = ~(layer_0[973] ^ layer_0[2515]); 
    assign out[1021] = ~layer_0[1977]; 
    assign out[1022] = layer_0[1580] ^ layer_0[1568]; 
    assign out[1023] = ~layer_0[211]; 
    assign out[1024] = ~(layer_0[1293] | layer_0[378]); 
    assign out[1025] = layer_0[356]; 
    assign out[1026] = layer_0[1162] & layer_0[21]; 
    assign out[1027] = ~(layer_0[1925] ^ layer_0[2140]); 
    assign out[1028] = layer_0[2406] & ~layer_0[1613]; 
    assign out[1029] = ~(layer_0[1034] ^ layer_0[607]); 
    assign out[1030] = layer_0[1735] & layer_0[1942]; 
    assign out[1031] = ~(layer_0[2271] | layer_0[1625]); 
    assign out[1032] = ~layer_0[494]; 
    assign out[1033] = ~layer_0[955]; 
    assign out[1034] = ~(layer_0[2436] | layer_0[1609]); 
    assign out[1035] = layer_0[1657] ^ layer_0[1898]; 
    assign out[1036] = ~layer_0[1797] | (layer_0[805] & layer_0[1797]); 
    assign out[1037] = layer_0[2231]; 
    assign out[1038] = ~layer_0[1228]; 
    assign out[1039] = layer_0[275]; 
    assign out[1040] = ~(layer_0[2064] ^ layer_0[198]); 
    assign out[1041] = ~layer_0[1649]; 
    assign out[1042] = ~layer_0[2532] | (layer_0[125] & layer_0[2532]); 
    assign out[1043] = layer_0[1087] ^ layer_0[1634]; 
    assign out[1044] = layer_0[360] ^ layer_0[844]; 
    assign out[1045] = layer_0[1668] & ~layer_0[252]; 
    assign out[1046] = ~layer_0[329]; 
    assign out[1047] = layer_0[2181] ^ layer_0[2163]; 
    assign out[1048] = ~layer_0[372]; 
    assign out[1049] = layer_0[1267]; 
    assign out[1050] = ~(layer_0[908] & layer_0[2018]); 
    assign out[1051] = layer_0[1656] & layer_0[457]; 
    assign out[1052] = layer_0[1074] | layer_0[1299]; 
    assign out[1053] = layer_0[852] ^ layer_0[1928]; 
    assign out[1054] = ~(layer_0[1537] ^ layer_0[902]); 
    assign out[1055] = layer_0[1192] & layer_0[1645]; 
    assign out[1056] = layer_0[1229] ^ layer_0[405]; 
    assign out[1057] = layer_0[354] | layer_0[2126]; 
    assign out[1058] = ~layer_0[2450]; 
    assign out[1059] = ~layer_0[1352]; 
    assign out[1060] = layer_0[233] & ~layer_0[2411]; 
    assign out[1061] = ~layer_0[1727]; 
    assign out[1062] = layer_0[240]; 
    assign out[1063] = ~(layer_0[1192] ^ layer_0[1013]); 
    assign out[1064] = ~(layer_0[985] ^ layer_0[658]); 
    assign out[1065] = ~(layer_0[1361] ^ layer_0[1883]); 
    assign out[1066] = ~layer_0[80] | (layer_0[89] & layer_0[80]); 
    assign out[1067] = layer_0[1120] ^ layer_0[1658]; 
    assign out[1068] = layer_0[1687]; 
    assign out[1069] = ~layer_0[1826] | (layer_0[1826] & layer_0[1036]); 
    assign out[1070] = ~layer_0[1185]; 
    assign out[1071] = layer_0[805]; 
    assign out[1072] = ~(layer_0[1504] ^ layer_0[1334]); 
    assign out[1073] = layer_0[1072]; 
    assign out[1074] = layer_0[62]; 
    assign out[1075] = ~layer_0[74]; 
    assign out[1076] = layer_0[1113]; 
    assign out[1077] = layer_0[2198]; 
    assign out[1078] = ~(layer_0[1662] | layer_0[1092]); 
    assign out[1079] = layer_0[847] & layer_0[1777]; 
    assign out[1080] = ~(layer_0[1426] ^ layer_0[72]); 
    assign out[1081] = ~(layer_0[2149] & layer_0[1908]); 
    assign out[1082] = layer_0[2263] & ~layer_0[2557]; 
    assign out[1083] = ~layer_0[2199] | (layer_0[2199] & layer_0[2124]); 
    assign out[1084] = ~layer_0[93]; 
    assign out[1085] = ~(layer_0[484] & layer_0[503]); 
    assign out[1086] = layer_0[21] & ~layer_0[794]; 
    assign out[1087] = layer_0[148] & ~layer_0[1609]; 
    assign out[1088] = layer_0[1274]; 
    assign out[1089] = layer_0[1395] & ~layer_0[215]; 
    assign out[1090] = ~(layer_0[699] ^ layer_0[77]); 
    assign out[1091] = ~layer_0[2459]; 
    assign out[1092] = layer_0[2263]; 
    assign out[1093] = ~layer_0[1188]; 
    assign out[1094] = layer_0[1444] & ~layer_0[918]; 
    assign out[1095] = ~layer_0[1188]; 
    assign out[1096] = ~layer_0[1793]; 
    assign out[1097] = layer_0[1424]; 
    assign out[1098] = layer_0[1314] & ~layer_0[1767]; 
    assign out[1099] = ~(layer_0[1664] ^ layer_0[1557]); 
    assign out[1100] = layer_0[2533] ^ layer_0[802]; 
    assign out[1101] = ~layer_0[2331]; 
    assign out[1102] = layer_0[1154]; 
    assign out[1103] = ~(layer_0[171] & layer_0[1983]); 
    assign out[1104] = ~layer_0[309]; 
    assign out[1105] = ~layer_0[83]; 
    assign out[1106] = layer_0[560] & ~layer_0[2212]; 
    assign out[1107] = ~(layer_0[884] | layer_0[2114]); 
    assign out[1108] = ~(layer_0[475] & layer_0[1170]); 
    assign out[1109] = layer_0[1094]; 
    assign out[1110] = ~layer_0[2256]; 
    assign out[1111] = ~(layer_0[1286] & layer_0[875]); 
    assign out[1112] = ~(layer_0[306] & layer_0[2163]); 
    assign out[1113] = ~layer_0[477]; 
    assign out[1114] = ~layer_0[93]; 
    assign out[1115] = ~layer_0[1047]; 
    assign out[1116] = layer_0[1134] & ~layer_0[1733]; 
    assign out[1117] = ~layer_0[813]; 
    assign out[1118] = layer_0[846] & ~layer_0[326]; 
    assign out[1119] = ~(layer_0[1957] | layer_0[1757]); 
    assign out[1120] = layer_0[637] ^ layer_0[392]; 
    assign out[1121] = ~(layer_0[471] & layer_0[2030]); 
    assign out[1122] = ~layer_0[158]; 
    assign out[1123] = layer_0[2296] ^ layer_0[519]; 
    assign out[1124] = ~layer_0[2363]; 
    assign out[1125] = layer_0[2046] & ~layer_0[1075]; 
    assign out[1126] = ~layer_0[469]; 
    assign out[1127] = ~layer_0[2092]; 
    assign out[1128] = ~layer_0[281]; 
    assign out[1129] = layer_0[924]; 
    assign out[1130] = ~layer_0[537] | (layer_0[537] & layer_0[55]); 
    assign out[1131] = ~(layer_0[558] ^ layer_0[1681]); 
    assign out[1132] = ~layer_0[137]; 
    assign out[1133] = ~(layer_0[952] ^ layer_0[1876]); 
    assign out[1134] = ~layer_0[1625]; 
    assign out[1135] = ~layer_0[1982] | (layer_0[1982] & layer_0[738]); 
    assign out[1136] = ~(layer_0[1665] ^ layer_0[833]); 
    assign out[1137] = layer_0[2065]; 
    assign out[1138] = layer_0[1596] & ~layer_0[1847]; 
    assign out[1139] = ~layer_0[535]; 
    assign out[1140] = ~layer_0[1927] | (layer_0[1927] & layer_0[71]); 
    assign out[1141] = layer_0[805] & layer_0[607]; 
    assign out[1142] = ~layer_0[2448] | (layer_0[2448] & layer_0[1329]); 
    assign out[1143] = ~(layer_0[1304] ^ layer_0[1229]); 
    assign out[1144] = ~(layer_0[1106] | layer_0[590]); 
    assign out[1145] = ~(layer_0[1538] ^ layer_0[559]); 
    assign out[1146] = ~(layer_0[308] | layer_0[2531]); 
    assign out[1147] = ~layer_0[946]; 
    assign out[1148] = layer_0[290]; 
    assign out[1149] = ~layer_0[58]; 
    assign out[1150] = layer_0[2526] ^ layer_0[7]; 
    assign out[1151] = ~(layer_0[741] & layer_0[2163]); 
    assign out[1152] = layer_0[388] & ~layer_0[559]; 
    assign out[1153] = ~(layer_0[2448] & layer_0[693]); 
    assign out[1154] = ~(layer_0[1222] ^ layer_0[2058]); 
    assign out[1155] = ~(layer_0[481] | layer_0[1982]); 
    assign out[1156] = layer_0[2218] ^ layer_0[1100]; 
    assign out[1157] = layer_0[2340] ^ layer_0[28]; 
    assign out[1158] = layer_0[1227]; 
    assign out[1159] = layer_0[1203] ^ layer_0[829]; 
    assign out[1160] = layer_0[2509] ^ layer_0[232]; 
    assign out[1161] = layer_0[1605] ^ layer_0[1676]; 
    assign out[1162] = layer_0[2414]; 
    assign out[1163] = ~(layer_0[741] ^ layer_0[322]); 
    assign out[1164] = layer_0[842] & ~layer_0[1561]; 
    assign out[1165] = ~(layer_0[136] & layer_0[1689]); 
    assign out[1166] = ~(layer_0[1030] ^ layer_0[1429]); 
    assign out[1167] = layer_0[1206] & layer_0[988]; 
    assign out[1168] = layer_0[778] ^ layer_0[712]; 
    assign out[1169] = ~(layer_0[2017] & layer_0[195]); 
    assign out[1170] = ~(layer_0[283] ^ layer_0[48]); 
    assign out[1171] = ~layer_0[1142] | (layer_0[1804] & layer_0[1142]); 
    assign out[1172] = ~(layer_0[2244] ^ layer_0[621]); 
    assign out[1173] = ~(layer_0[1444] ^ layer_0[1001]); 
    assign out[1174] = layer_0[1676]; 
    assign out[1175] = ~layer_0[929] | (layer_0[1043] & layer_0[929]); 
    assign out[1176] = layer_0[2228] & ~layer_0[1865]; 
    assign out[1177] = layer_0[1151] ^ layer_0[1486]; 
    assign out[1178] = layer_0[1481]; 
    assign out[1179] = layer_0[1831] & ~layer_0[460]; 
    assign out[1180] = layer_0[1430] ^ layer_0[2396]; 
    assign out[1181] = ~(layer_0[412] ^ layer_0[1916]); 
    assign out[1182] = layer_0[1168]; 
    assign out[1183] = layer_0[454] & layer_0[1103]; 
    assign out[1184] = ~(layer_0[1326] | layer_0[1038]); 
    assign out[1185] = ~(layer_0[1363] | layer_0[136]); 
    assign out[1186] = ~(layer_0[1244] ^ layer_0[425]); 
    assign out[1187] = ~(layer_0[1936] | layer_0[85]); 
    assign out[1188] = layer_0[1475]; 
    assign out[1189] = ~layer_0[1684]; 
    assign out[1190] = ~layer_0[2469]; 
    assign out[1191] = layer_0[1034] & ~layer_0[1328]; 
    assign out[1192] = ~(layer_0[49] | layer_0[167]); 
    assign out[1193] = layer_0[2382] ^ layer_0[2079]; 
    assign out[1194] = layer_0[373] ^ layer_0[1225]; 
    assign out[1195] = layer_0[1162] & ~layer_0[4]; 
    assign out[1196] = ~layer_0[137]; 
    assign out[1197] = ~(layer_0[335] | layer_0[2061]); 
    assign out[1198] = layer_0[2389]; 
    assign out[1199] = layer_0[2040] & layer_0[1162]; 
    assign out[1200] = ~layer_0[884]; 
    assign out[1201] = ~(layer_0[1657] & layer_0[1303]); 
    assign out[1202] = ~(layer_0[16] ^ layer_0[454]); 
    assign out[1203] = layer_0[2105] & layer_0[153]; 
    assign out[1204] = layer_0[1488]; 
    assign out[1205] = layer_0[515]; 
    assign out[1206] = layer_0[2414]; 
    assign out[1207] = ~(layer_0[218] ^ layer_0[683]); 
    assign out[1208] = ~layer_0[1631]; 
    assign out[1209] = layer_0[959] & ~layer_0[940]; 
    assign out[1210] = ~(layer_0[28] & layer_0[581]); 
    assign out[1211] = layer_0[764]; 
    assign out[1212] = ~layer_0[2427]; 
    assign out[1213] = layer_0[608] | layer_0[750]; 
    assign out[1214] = layer_0[1006]; 
    assign out[1215] = layer_0[1833] & ~layer_0[2150]; 
    assign out[1216] = layer_0[101] ^ layer_0[2444]; 
    assign out[1217] = ~(layer_0[1057] | layer_0[395]); 
    assign out[1218] = ~(layer_0[2340] ^ layer_0[838]); 
    assign out[1219] = layer_0[2068]; 
    assign out[1220] = layer_0[10] & ~layer_0[2378]; 
    assign out[1221] = ~(layer_0[1813] ^ layer_0[2241]); 
    assign out[1222] = layer_0[1405]; 
    assign out[1223] = ~(layer_0[2256] | layer_0[2402]); 
    assign out[1224] = ~layer_0[93] | (layer_0[93] & layer_0[657]); 
    assign out[1225] = ~layer_0[2230] | (layer_0[2230] & layer_0[1393]); 
    assign out[1226] = layer_0[1829] & ~layer_0[1982]; 
    assign out[1227] = layer_0[959]; 
    assign out[1228] = ~layer_0[1556]; 
    assign out[1229] = ~layer_0[1296]; 
    assign out[1230] = ~(layer_0[1652] & layer_0[1927]); 
    assign out[1231] = layer_0[2508]; 
    assign out[1232] = ~(layer_0[184] | layer_0[1235]); 
    assign out[1233] = ~(layer_0[2505] ^ layer_0[969]); 
    assign out[1234] = ~layer_0[1260]; 
    assign out[1235] = ~(layer_0[598] | layer_0[4]); 
    assign out[1236] = ~layer_0[357] | (layer_0[2213] & layer_0[357]); 
    assign out[1237] = ~(layer_0[1259] | layer_0[206]); 
    assign out[1238] = layer_0[357] ^ layer_0[785]; 
    assign out[1239] = layer_0[1788]; 
    assign out[1240] = layer_0[2484]; 
    assign out[1241] = layer_0[520]; 
    assign out[1242] = layer_0[2514] ^ layer_0[2393]; 
    assign out[1243] = layer_0[431]; 
    assign out[1244] = ~(layer_0[1026] | layer_0[1463]); 
    assign out[1245] = ~layer_0[455] | (layer_0[455] & layer_0[873]); 
    assign out[1246] = ~layer_0[587] | (layer_0[587] & layer_0[291]); 
    assign out[1247] = layer_0[170] ^ layer_0[649]; 
    assign out[1248] = ~(layer_0[1005] ^ layer_0[2126]); 
    assign out[1249] = ~layer_0[2033]; 
    assign out[1250] = layer_0[193] & ~layer_0[1204]; 
    assign out[1251] = layer_0[2004] & layer_0[591]; 
    assign out[1252] = ~(layer_0[1980] ^ layer_0[2011]); 
    assign out[1253] = ~(layer_0[1652] | layer_0[770]); 
    assign out[1254] = layer_0[125] & ~layer_0[115]; 
    assign out[1255] = layer_0[2097] & ~layer_0[2312]; 
    assign out[1256] = layer_0[700]; 
    assign out[1257] = layer_0[1246]; 
    assign out[1258] = ~layer_0[1941]; 
    assign out[1259] = ~layer_0[544]; 
    assign out[1260] = layer_0[197]; 
    assign out[1261] = layer_0[2014] & layer_0[2190]; 
    assign out[1262] = ~(layer_0[2483] ^ layer_0[2291]); 
    assign out[1263] = ~layer_0[439]; 
    assign out[1264] = ~layer_0[1185]; 
    assign out[1265] = layer_0[1498]; 
    assign out[1266] = layer_0[2311] ^ layer_0[1078]; 
    assign out[1267] = layer_0[2059] ^ layer_0[1340]; 
    assign out[1268] = layer_0[1782] ^ layer_0[658]; 
    assign out[1269] = ~layer_0[144]; 
    assign out[1270] = layer_0[1889]; 
    assign out[1271] = layer_0[1165] | layer_0[1894]; 
    assign out[1272] = layer_0[1761] & layer_0[1942]; 
    assign out[1273] = ~layer_0[1484]; 
    assign out[1274] = layer_0[2383] ^ layer_0[2554]; 
    assign out[1275] = ~(layer_0[1053] ^ layer_0[1362]); 
    assign out[1276] = layer_0[385]; 
    assign out[1277] = ~(layer_0[784] ^ layer_0[1221]); 
    assign out[1278] = ~(layer_0[2442] ^ layer_0[2090]); 
    assign out[1279] = ~layer_0[2004]; 
    assign out[1280] = ~(layer_0[508] ^ layer_0[1190]); 
    assign out[1281] = layer_0[543] ^ layer_0[1765]; 
    assign out[1282] = layer_0[2501]; 
    assign out[1283] = layer_0[1317]; 
    assign out[1284] = layer_0[434]; 
    assign out[1285] = ~(layer_0[384] ^ layer_0[1284]); 
    assign out[1286] = ~(layer_0[691] ^ layer_0[10]); 
    assign out[1287] = ~(layer_0[339] ^ layer_0[1993]); 
    assign out[1288] = ~(layer_0[538] & layer_0[706]); 
    assign out[1289] = ~(layer_0[2505] ^ layer_0[2061]); 
    assign out[1290] = layer_0[1403] & ~layer_0[1628]; 
    assign out[1291] = ~(layer_0[1748] ^ layer_0[973]); 
    assign out[1292] = layer_0[602] ^ layer_0[777]; 
    assign out[1293] = layer_0[1005] ^ layer_0[826]; 
    assign out[1294] = ~(layer_0[1579] ^ layer_0[1833]); 
    assign out[1295] = ~layer_0[2449]; 
    assign out[1296] = ~layer_0[1043]; 
    assign out[1297] = layer_0[402]; 
    assign out[1298] = layer_0[2080] | layer_0[856]; 
    assign out[1299] = layer_0[1766] | layer_0[1612]; 
    assign out[1300] = layer_0[1878] ^ layer_0[1127]; 
    assign out[1301] = ~(layer_0[1510] ^ layer_0[664]); 
    assign out[1302] = ~(layer_0[219] ^ layer_0[2182]); 
    assign out[1303] = ~(layer_0[2356] ^ layer_0[877]); 
    assign out[1304] = layer_0[2232] ^ layer_0[2160]; 
    assign out[1305] = layer_0[2256] | layer_0[1849]; 
    assign out[1306] = layer_0[229]; 
    assign out[1307] = ~layer_0[1959]; 
    assign out[1308] = ~layer_0[414]; 
    assign out[1309] = ~(layer_0[339] | layer_0[2384]); 
    assign out[1310] = ~(layer_0[1369] ^ layer_0[18]); 
    assign out[1311] = layer_0[640] & ~layer_0[901]; 
    assign out[1312] = ~(layer_0[2550] ^ layer_0[1512]); 
    assign out[1313] = layer_0[1783] ^ layer_0[283]; 
    assign out[1314] = layer_0[11] | layer_0[267]; 
    assign out[1315] = layer_0[1173] ^ layer_0[2000]; 
    assign out[1316] = ~(layer_0[1607] | layer_0[2048]); 
    assign out[1317] = ~layer_0[2332]; 
    assign out[1318] = ~layer_0[396]; 
    assign out[1319] = layer_0[1010]; 
    assign out[1320] = layer_0[2418] ^ layer_0[1107]; 
    assign out[1321] = layer_0[35] ^ layer_0[1780]; 
    assign out[1322] = layer_0[109]; 
    assign out[1323] = layer_0[1334]; 
    assign out[1324] = layer_0[1442] ^ layer_0[1189]; 
    assign out[1325] = ~(layer_0[192] ^ layer_0[2544]); 
    assign out[1326] = ~(layer_0[356] ^ layer_0[1918]); 
    assign out[1327] = ~(layer_0[2379] ^ layer_0[1382]); 
    assign out[1328] = layer_0[2102] ^ layer_0[2042]; 
    assign out[1329] = layer_0[1777] & ~layer_0[677]; 
    assign out[1330] = ~(layer_0[2486] ^ layer_0[972]); 
    assign out[1331] = ~layer_0[10]; 
    assign out[1332] = ~(layer_0[1023] ^ layer_0[114]); 
    assign out[1333] = layer_0[1366] & ~layer_0[1338]; 
    assign out[1334] = layer_0[726]; 
    assign out[1335] = ~layer_0[1176]; 
    assign out[1336] = ~layer_0[1271]; 
    assign out[1337] = layer_0[424] & ~layer_0[1338]; 
    assign out[1338] = ~layer_0[2081]; 
    assign out[1339] = ~layer_0[2505]; 
    assign out[1340] = ~layer_0[2052] | (layer_0[2052] & layer_0[1604]); 
    assign out[1341] = layer_0[1833] ^ layer_0[117]; 
    assign out[1342] = layer_0[1387]; 
    assign out[1343] = layer_0[1793] & layer_0[875]; 
    assign out[1344] = ~layer_0[599]; 
    assign out[1345] = ~(layer_0[1404] ^ layer_0[462]); 
    assign out[1346] = ~(layer_0[2365] ^ layer_0[1717]); 
    assign out[1347] = ~layer_0[1418] | (layer_0[1418] & layer_0[1367]); 
    assign out[1348] = layer_0[2031]; 
    assign out[1349] = layer_0[1832]; 
    assign out[1350] = ~layer_0[1375] | (layer_0[1375] & layer_0[2541]); 
    assign out[1351] = ~layer_0[848] | (layer_0[848] & layer_0[836]); 
    assign out[1352] = ~layer_0[548]; 
    assign out[1353] = ~(layer_0[227] ^ layer_0[357]); 
    assign out[1354] = ~(layer_0[670] ^ layer_0[728]); 
    assign out[1355] = layer_0[1832]; 
    assign out[1356] = layer_0[127]; 
    assign out[1357] = layer_0[2240]; 
    assign out[1358] = ~(layer_0[1140] & layer_0[581]); 
    assign out[1359] = ~layer_0[1632] | (layer_0[260] & layer_0[1632]); 
    assign out[1360] = layer_0[921] & ~layer_0[912]; 
    assign out[1361] = layer_0[424] | layer_0[435]; 
    assign out[1362] = layer_0[2385] & layer_0[2541]; 
    assign out[1363] = layer_0[173] & ~layer_0[1643]; 
    assign out[1364] = ~(layer_0[198] & layer_0[98]); 
    assign out[1365] = layer_0[1276]; 
    assign out[1366] = ~(layer_0[2229] ^ layer_0[1558]); 
    assign out[1367] = layer_0[1226]; 
    assign out[1368] = layer_0[2443] | layer_0[137]; 
    assign out[1369] = layer_0[2176]; 
    assign out[1370] = layer_0[1938] & ~layer_0[1141]; 
    assign out[1371] = layer_0[1613] ^ layer_0[275]; 
    assign out[1372] = ~(layer_0[1726] | layer_0[423]); 
    assign out[1373] = layer_0[1233] & ~layer_0[2336]; 
    assign out[1374] = ~layer_0[2005]; 
    assign out[1375] = layer_0[114] & ~layer_0[1807]; 
    assign out[1376] = ~layer_0[426] | (layer_0[2466] & layer_0[426]); 
    assign out[1377] = ~layer_0[1132]; 
    assign out[1378] = layer_0[1968]; 
    assign out[1379] = layer_0[2292] ^ layer_0[1178]; 
    assign out[1380] = ~layer_0[1435]; 
    assign out[1381] = ~layer_0[917]; 
    assign out[1382] = layer_0[434] ^ layer_0[530]; 
    assign out[1383] = ~layer_0[1770] | (layer_0[1770] & layer_0[1981]); 
    assign out[1384] = ~(layer_0[1628] | layer_0[2279]); 
    assign out[1385] = ~(layer_0[1054] & layer_0[1154]); 
    assign out[1386] = layer_0[1291]; 
    assign out[1387] = ~(layer_0[1534] ^ layer_0[1842]); 
    assign out[1388] = ~layer_0[2431]; 
    assign out[1389] = layer_0[1252]; 
    assign out[1390] = layer_0[305] & layer_0[113]; 
    assign out[1391] = layer_0[511] ^ layer_0[707]; 
    assign out[1392] = ~(layer_0[1988] ^ layer_0[555]); 
    assign out[1393] = layer_0[1051] ^ layer_0[279]; 
    assign out[1394] = ~(layer_0[401] ^ layer_0[2556]); 
    assign out[1395] = ~layer_0[651]; 
    assign out[1396] = ~layer_0[20]; 
    assign out[1397] = ~layer_0[1629]; 
    assign out[1398] = layer_0[863] ^ layer_0[135]; 
    assign out[1399] = layer_0[2330] ^ layer_0[1599]; 
    assign out[1400] = ~layer_0[1382] | (layer_0[1382] & layer_0[531]); 
    assign out[1401] = ~layer_0[1779]; 
    assign out[1402] = ~(layer_0[222] ^ layer_0[61]); 
    assign out[1403] = ~layer_0[1108]; 
    assign out[1404] = ~(layer_0[2395] ^ layer_0[498]); 
    assign out[1405] = layer_0[721] & ~layer_0[426]; 
    assign out[1406] = ~layer_0[759] | (layer_0[424] & layer_0[759]); 
    assign out[1407] = layer_0[1509] & ~layer_0[1588]; 
    assign out[1408] = ~(layer_0[1271] | layer_0[1583]); 
    assign out[1409] = ~(layer_0[2513] ^ layer_0[1730]); 
    assign out[1410] = layer_0[640] & layer_0[1459]; 
    assign out[1411] = layer_0[854]; 
    assign out[1412] = layer_0[1793] | layer_0[1305]; 
    assign out[1413] = ~layer_0[35] | (layer_0[847] & layer_0[35]); 
    assign out[1414] = layer_0[329]; 
    assign out[1415] = layer_0[361] & ~layer_0[1623]; 
    assign out[1416] = ~(layer_0[1667] ^ layer_0[451]); 
    assign out[1417] = ~layer_0[1619] | (layer_0[14] & layer_0[1619]); 
    assign out[1418] = ~(layer_0[1654] ^ layer_0[2425]); 
    assign out[1419] = layer_0[837]; 
    assign out[1420] = layer_0[1387]; 
    assign out[1421] = layer_0[1219] ^ layer_0[1084]; 
    assign out[1422] = ~layer_0[1607]; 
    assign out[1423] = layer_0[2089]; 
    assign out[1424] = layer_0[196] | layer_0[1233]; 
    assign out[1425] = layer_0[547]; 
    assign out[1426] = ~layer_0[712]; 
    assign out[1427] = ~(layer_0[2431] | layer_0[881]); 
    assign out[1428] = ~(layer_0[1070] ^ layer_0[2411]); 
    assign out[1429] = layer_0[2330] ^ layer_0[2434]; 
    assign out[1430] = layer_0[1183]; 
    assign out[1431] = layer_0[2307] ^ layer_0[912]; 
    assign out[1432] = ~layer_0[1135] | (layer_0[1135] & layer_0[1358]); 
    assign out[1433] = ~(layer_0[970] & layer_0[41]); 
    assign out[1434] = layer_0[1014] ^ layer_0[1786]; 
    assign out[1435] = layer_0[593]; 
    assign out[1436] = layer_0[2352] ^ layer_0[1035]; 
    assign out[1437] = layer_0[574]; 
    assign out[1438] = layer_0[2260]; 
    assign out[1439] = layer_0[420] ^ layer_0[1623]; 
    assign out[1440] = ~layer_0[2384]; 
    assign out[1441] = layer_0[875]; 
    assign out[1442] = ~layer_0[1816]; 
    assign out[1443] = ~(layer_0[216] ^ layer_0[2315]); 
    assign out[1444] = ~(layer_0[1987] ^ layer_0[2133]); 
    assign out[1445] = ~layer_0[1534] | (layer_0[1534] & layer_0[542]); 
    assign out[1446] = layer_0[795]; 
    assign out[1447] = layer_0[1222]; 
    assign out[1448] = layer_0[2466] & layer_0[2210]; 
    assign out[1449] = layer_0[586] | layer_0[259]; 
    assign out[1450] = ~(layer_0[761] & layer_0[1882]); 
    assign out[1451] = layer_0[1256]; 
    assign out[1452] = layer_0[534] & layer_0[858]; 
    assign out[1453] = layer_0[1466] ^ layer_0[1182]; 
    assign out[1454] = ~layer_0[2086]; 
    assign out[1455] = layer_0[2298]; 
    assign out[1456] = layer_0[646]; 
    assign out[1457] = ~(layer_0[11] ^ layer_0[2034]); 
    assign out[1458] = layer_0[2123] ^ layer_0[2316]; 
    assign out[1459] = ~(layer_0[1693] ^ layer_0[1307]); 
    assign out[1460] = ~layer_0[2111]; 
    assign out[1461] = layer_0[375] ^ layer_0[1410]; 
    assign out[1462] = layer_0[1427] | layer_0[2551]; 
    assign out[1463] = ~(layer_0[870] ^ layer_0[756]); 
    assign out[1464] = ~layer_0[712]; 
    assign out[1465] = layer_0[2130]; 
    assign out[1466] = ~(layer_0[561] ^ layer_0[218]); 
    assign out[1467] = ~(layer_0[835] ^ layer_0[605]); 
    assign out[1468] = layer_0[1878] ^ layer_0[1449]; 
    assign out[1469] = ~layer_0[1599]; 
    assign out[1470] = layer_0[1441] ^ layer_0[151]; 
    assign out[1471] = ~(layer_0[1961] ^ layer_0[1006]); 
    assign out[1472] = ~(layer_0[58] ^ layer_0[483]); 
    assign out[1473] = ~layer_0[684] | (layer_0[2465] & layer_0[684]); 
    assign out[1474] = layer_0[2044] ^ layer_0[14]; 
    assign out[1475] = layer_0[2462] & ~layer_0[1668]; 
    assign out[1476] = ~(layer_0[1036] | layer_0[665]); 
    assign out[1477] = layer_0[137]; 
    assign out[1478] = ~(layer_0[811] ^ layer_0[337]); 
    assign out[1479] = ~layer_0[234]; 
    assign out[1480] = ~(layer_0[458] | layer_0[1457]); 
    assign out[1481] = ~layer_0[64]; 
    assign out[1482] = ~(layer_0[513] | layer_0[1372]); 
    assign out[1483] = ~(layer_0[765] & layer_0[143]); 
    assign out[1484] = ~layer_0[1407]; 
    assign out[1485] = layer_0[870]; 
    assign out[1486] = layer_0[2538] | layer_0[1301]; 
    assign out[1487] = layer_0[536] ^ layer_0[977]; 
    assign out[1488] = layer_0[2190] ^ layer_0[915]; 
    assign out[1489] = ~layer_0[1779] | (layer_0[1779] & layer_0[534]); 
    assign out[1490] = layer_0[533] ^ layer_0[303]; 
    assign out[1491] = ~layer_0[490]; 
    assign out[1492] = layer_0[1465] ^ layer_0[1707]; 
    assign out[1493] = layer_0[2466]; 
    assign out[1494] = layer_0[2473] & layer_0[1612]; 
    assign out[1495] = ~(layer_0[2326] ^ layer_0[1173]); 
    assign out[1496] = ~(layer_0[2316] | layer_0[1672]); 
    assign out[1497] = ~layer_0[1478]; 
    assign out[1498] = layer_0[605] ^ layer_0[1789]; 
    assign out[1499] = layer_0[2435] | layer_0[1275]; 
    assign out[1500] = layer_0[1097]; 
    assign out[1501] = ~layer_0[2468] | (layer_0[2468] & layer_0[2260]); 
    assign out[1502] = ~(layer_0[908] ^ layer_0[1638]); 
    assign out[1503] = layer_0[386]; 
    assign out[1504] = ~layer_0[570]; 
    assign out[1505] = layer_0[1502]; 
    assign out[1506] = layer_0[229] | layer_0[1189]; 
    assign out[1507] = layer_0[1212]; 
    assign out[1508] = layer_0[280]; 
    assign out[1509] = ~layer_0[2255] | (layer_0[2255] & layer_0[1517]); 
    assign out[1510] = layer_0[1252]; 
    assign out[1511] = ~(layer_0[197] | layer_0[1372]); 
    assign out[1512] = layer_0[122]; 
    assign out[1513] = layer_0[2209] & ~layer_0[754]; 
    assign out[1514] = layer_0[2324] & layer_0[670]; 
    assign out[1515] = ~layer_0[377]; 
    assign out[1516] = layer_0[409]; 
    assign out[1517] = layer_0[330] ^ layer_0[39]; 
    assign out[1518] = ~(layer_0[108] ^ layer_0[1385]); 
    assign out[1519] = ~(layer_0[2440] ^ layer_0[2400]); 
    assign out[1520] = ~(layer_0[1528] ^ layer_0[1972]); 
    assign out[1521] = layer_0[23] & layer_0[1755]; 
    assign out[1522] = ~layer_0[1629]; 
    assign out[1523] = ~(layer_0[2422] ^ layer_0[661]); 
    assign out[1524] = layer_0[1317]; 
    assign out[1525] = layer_0[409] ^ layer_0[769]; 
    assign out[1526] = layer_0[1165] ^ layer_0[2422]; 
    assign out[1527] = ~layer_0[706] | (layer_0[799] & layer_0[706]); 
    assign out[1528] = ~layer_0[562] | (layer_0[2335] & layer_0[562]); 
    assign out[1529] = layer_0[835] & ~layer_0[432]; 
    assign out[1530] = layer_0[2031] & ~layer_0[519]; 
    assign out[1531] = layer_0[2244]; 
    assign out[1532] = layer_0[2539] & ~layer_0[90]; 
    assign out[1533] = ~layer_0[237] | (layer_0[79] & layer_0[237]); 
    assign out[1534] = ~(layer_0[2315] | layer_0[1813]); 
    assign out[1535] = ~layer_0[1501] | (layer_0[1501] & layer_0[2296]); 
    assign out[1536] = ~layer_0[250]; 
    assign out[1537] = ~layer_0[525] | (layer_0[655] & layer_0[525]); 
    assign out[1538] = ~(layer_0[1001] & layer_0[1863]); 
    assign out[1539] = layer_0[2004]; 
    assign out[1540] = layer_0[397] ^ layer_0[2109]; 
    assign out[1541] = layer_0[1352] & ~layer_0[2373]; 
    assign out[1542] = ~(layer_0[1545] | layer_0[82]); 
    assign out[1543] = layer_0[811] ^ layer_0[166]; 
    assign out[1544] = layer_0[368] ^ layer_0[2015]; 
    assign out[1545] = ~(layer_0[2334] ^ layer_0[7]); 
    assign out[1546] = ~layer_0[2401]; 
    assign out[1547] = ~layer_0[1262]; 
    assign out[1548] = layer_0[942]; 
    assign out[1549] = ~(layer_0[57] | layer_0[523]); 
    assign out[1550] = ~layer_0[2177] | (layer_0[1440] & layer_0[2177]); 
    assign out[1551] = layer_0[1988] & ~layer_0[2446]; 
    assign out[1552] = ~layer_0[2299]; 
    assign out[1553] = ~(layer_0[2314] | layer_0[421]); 
    assign out[1554] = ~(layer_0[940] | layer_0[871]); 
    assign out[1555] = ~layer_0[2484]; 
    assign out[1556] = layer_0[313] & ~layer_0[1208]; 
    assign out[1557] = ~(layer_0[1062] ^ layer_0[2294]); 
    assign out[1558] = layer_0[1759]; 
    assign out[1559] = ~(layer_0[49] ^ layer_0[2269]); 
    assign out[1560] = ~layer_0[469]; 
    assign out[1561] = ~layer_0[1484]; 
    assign out[1562] = layer_0[1171] & ~layer_0[1429]; 
    assign out[1563] = layer_0[1636]; 
    assign out[1564] = layer_0[165] | layer_0[922]; 
    assign out[1565] = ~(layer_0[1762] | layer_0[1310]); 
    assign out[1566] = ~(layer_0[108] ^ layer_0[663]); 
    assign out[1567] = layer_0[1570] & ~layer_0[1452]; 
    assign out[1568] = ~layer_0[1]; 
    assign out[1569] = layer_0[2106]; 
    assign out[1570] = layer_0[437] & ~layer_0[1657]; 
    assign out[1571] = layer_0[2493]; 
    assign out[1572] = layer_0[2546] | layer_0[1096]; 
    assign out[1573] = layer_0[2558] | layer_0[1136]; 
    assign out[1574] = layer_0[603] & layer_0[1184]; 
    assign out[1575] = layer_0[1846]; 
    assign out[1576] = layer_0[354]; 
    assign out[1577] = ~(layer_0[1863] | layer_0[573]); 
    assign out[1578] = ~(layer_0[498] ^ layer_0[2082]); 
    assign out[1579] = ~(layer_0[2517] | layer_0[697]); 
    assign out[1580] = layer_0[1520]; 
    assign out[1581] = layer_0[2071]; 
    assign out[1582] = ~layer_0[573]; 
    assign out[1583] = layer_0[526] | layer_0[423]; 
    assign out[1584] = layer_0[1367] & layer_0[335]; 
    assign out[1585] = ~(layer_0[788] | layer_0[2314]); 
    assign out[1586] = layer_0[379] ^ layer_0[1854]; 
    assign out[1587] = layer_0[143] & ~layer_0[1075]; 
    assign out[1588] = layer_0[897] & layer_0[2319]; 
    assign out[1589] = ~(layer_0[101] & layer_0[1175]); 
    assign out[1590] = ~(layer_0[222] | layer_0[2277]); 
    assign out[1591] = ~layer_0[2007]; 
    assign out[1592] = layer_0[1759] & ~layer_0[1349]; 
    assign out[1593] = ~(layer_0[756] ^ layer_0[743]); 
    assign out[1594] = layer_0[409]; 
    assign out[1595] = ~layer_0[52]; 
    assign out[1596] = ~layer_0[2344]; 
    assign out[1597] = layer_0[1619]; 
    assign out[1598] = layer_0[1528]; 
    assign out[1599] = layer_0[1800] ^ layer_0[1977]; 
    assign out[1600] = ~layer_0[474]; 
    assign out[1601] = ~layer_0[368]; 
    assign out[1602] = layer_0[2070]; 
    assign out[1603] = ~layer_0[2379] | (layer_0[2379] & layer_0[560]); 
    assign out[1604] = ~layer_0[1166]; 
    assign out[1605] = layer_0[748]; 
    assign out[1606] = ~layer_0[2163]; 
    assign out[1607] = ~(layer_0[1834] ^ layer_0[2061]); 
    assign out[1608] = ~(layer_0[958] | layer_0[2481]); 
    assign out[1609] = layer_0[2489] & ~layer_0[241]; 
    assign out[1610] = layer_0[1530]; 
    assign out[1611] = layer_0[746] ^ layer_0[38]; 
    assign out[1612] = ~layer_0[2243]; 
    assign out[1613] = layer_0[551]; 
    assign out[1614] = ~layer_0[1879]; 
    assign out[1615] = layer_0[335]; 
    assign out[1616] = layer_0[1227]; 
    assign out[1617] = layer_0[2504] & ~layer_0[345]; 
    assign out[1618] = ~(layer_0[1506] | layer_0[1468]); 
    assign out[1619] = layer_0[2078] & ~layer_0[1065]; 
    assign out[1620] = ~layer_0[601]; 
    assign out[1621] = layer_0[2124] ^ layer_0[146]; 
    assign out[1622] = layer_0[913] & ~layer_0[510]; 
    assign out[1623] = ~(layer_0[762] ^ layer_0[1716]); 
    assign out[1624] = layer_0[932] & ~layer_0[1674]; 
    assign out[1625] = ~layer_0[759]; 
    assign out[1626] = layer_0[1454] & layer_0[412]; 
    assign out[1627] = ~layer_0[190]; 
    assign out[1628] = layer_0[2356] & layer_0[54]; 
    assign out[1629] = ~(layer_0[2497] ^ layer_0[1379]); 
    assign out[1630] = layer_0[1603] & ~layer_0[157]; 
    assign out[1631] = layer_0[932]; 
    assign out[1632] = layer_0[2347]; 
    assign out[1633] = layer_0[156]; 
    assign out[1634] = ~(layer_0[108] | layer_0[956]); 
    assign out[1635] = layer_0[2275]; 
    assign out[1636] = layer_0[1572] ^ layer_0[2088]; 
    assign out[1637] = layer_0[2055] & ~layer_0[1277]; 
    assign out[1638] = ~(layer_0[1436] | layer_0[46]); 
    assign out[1639] = ~(layer_0[515] ^ layer_0[86]); 
    assign out[1640] = layer_0[399] & ~layer_0[1093]; 
    assign out[1641] = ~(layer_0[2050] ^ layer_0[1145]); 
    assign out[1642] = ~layer_0[1310]; 
    assign out[1643] = ~(layer_0[1457] | layer_0[1226]); 
    assign out[1644] = ~(layer_0[559] | layer_0[2343]); 
    assign out[1645] = layer_0[1523] ^ layer_0[1965]; 
    assign out[1646] = ~layer_0[2177]; 
    assign out[1647] = ~(layer_0[102] & layer_0[1931]); 
    assign out[1648] = layer_0[126]; 
    assign out[1649] = layer_0[1559] ^ layer_0[1344]; 
    assign out[1650] = ~layer_0[605] | (layer_0[605] & layer_0[1477]); 
    assign out[1651] = layer_0[2237]; 
    assign out[1652] = ~layer_0[1982]; 
    assign out[1653] = ~(layer_0[2447] ^ layer_0[629]); 
    assign out[1654] = layer_0[2391]; 
    assign out[1655] = layer_0[1892] & layer_0[528]; 
    assign out[1656] = layer_0[2312]; 
    assign out[1657] = layer_0[1597]; 
    assign out[1658] = layer_0[1292] & ~layer_0[1185]; 
    assign out[1659] = ~(layer_0[1340] & layer_0[1279]); 
    assign out[1660] = layer_0[908] & ~layer_0[256]; 
    assign out[1661] = ~(layer_0[1210] ^ layer_0[1688]); 
    assign out[1662] = layer_0[1871] & ~layer_0[1495]; 
    assign out[1663] = ~layer_0[2026]; 
    assign out[1664] = layer_0[566]; 
    assign out[1665] = layer_0[1243]; 
    assign out[1666] = ~layer_0[247]; 
    assign out[1667] = layer_0[2144] ^ layer_0[1238]; 
    assign out[1668] = ~(layer_0[2551] | layer_0[1766]); 
    assign out[1669] = ~layer_0[2531]; 
    assign out[1670] = ~(layer_0[2422] | layer_0[2155]); 
    assign out[1671] = ~(layer_0[329] ^ layer_0[1903]); 
    assign out[1672] = ~layer_0[1202]; 
    assign out[1673] = ~(layer_0[1355] | layer_0[396]); 
    assign out[1674] = ~layer_0[1380] | (layer_0[1380] & layer_0[685]); 
    assign out[1675] = layer_0[897]; 
    assign out[1676] = ~(layer_0[77] & layer_0[2316]); 
    assign out[1677] = layer_0[224] & ~layer_0[2166]; 
    assign out[1678] = ~(layer_0[1768] ^ layer_0[1011]); 
    assign out[1679] = layer_0[86] & ~layer_0[795]; 
    assign out[1680] = ~(layer_0[1532] & layer_0[1937]); 
    assign out[1681] = layer_0[1907] ^ layer_0[1626]; 
    assign out[1682] = ~layer_0[712]; 
    assign out[1683] = layer_0[261] & layer_0[705]; 
    assign out[1684] = ~(layer_0[289] ^ layer_0[1027]); 
    assign out[1685] = ~layer_0[984]; 
    assign out[1686] = ~layer_0[1834] | (layer_0[548] & layer_0[1834]); 
    assign out[1687] = layer_0[1240] & ~layer_0[1903]; 
    assign out[1688] = layer_0[2216] & ~layer_0[689]; 
    assign out[1689] = layer_0[1802] ^ layer_0[1754]; 
    assign out[1690] = ~(layer_0[436] ^ layer_0[2357]); 
    assign out[1691] = layer_0[1988]; 
    assign out[1692] = layer_0[531] & ~layer_0[1774]; 
    assign out[1693] = layer_0[240] ^ layer_0[1878]; 
    assign out[1694] = layer_0[875] & ~layer_0[2236]; 
    assign out[1695] = layer_0[446]; 
    assign out[1696] = layer_0[611] & ~layer_0[2407]; 
    assign out[1697] = ~(layer_0[47] ^ layer_0[1552]); 
    assign out[1698] = layer_0[2036] ^ layer_0[1542]; 
    assign out[1699] = ~(layer_0[1419] ^ layer_0[2187]); 
    assign out[1700] = ~(layer_0[2404] ^ layer_0[58]); 
    assign out[1701] = layer_0[1136] ^ layer_0[622]; 
    assign out[1702] = ~layer_0[1562]; 
    assign out[1703] = layer_0[935]; 
    assign out[1704] = layer_0[2546] & layer_0[1782]; 
    assign out[1705] = layer_0[2038]; 
    assign out[1706] = layer_0[961] & layer_0[1177]; 
    assign out[1707] = ~(layer_0[1852] ^ layer_0[1395]); 
    assign out[1708] = ~layer_0[646]; 
    assign out[1709] = layer_0[2229] ^ layer_0[194]; 
    assign out[1710] = ~layer_0[524] | (layer_0[1655] & layer_0[524]); 
    assign out[1711] = ~(layer_0[1471] ^ layer_0[774]); 
    assign out[1712] = layer_0[1238] & ~layer_0[1186]; 
    assign out[1713] = layer_0[509] & ~layer_0[1525]; 
    assign out[1714] = ~(layer_0[2442] | layer_0[222]); 
    assign out[1715] = ~(layer_0[390] | layer_0[865]); 
    assign out[1716] = ~layer_0[193]; 
    assign out[1717] = layer_0[1878] ^ layer_0[2364]; 
    assign out[1718] = ~(layer_0[759] & layer_0[675]); 
    assign out[1719] = ~layer_0[188] | (layer_0[2309] & layer_0[188]); 
    assign out[1720] = ~layer_0[1774]; 
    assign out[1721] = layer_0[1096] & ~layer_0[1968]; 
    assign out[1722] = ~(layer_0[2048] ^ layer_0[1362]); 
    assign out[1723] = layer_0[2300] & layer_0[1304]; 
    assign out[1724] = layer_0[1995] & ~layer_0[2407]; 
    assign out[1725] = ~layer_0[2453]; 
    assign out[1726] = ~layer_0[1126] | (layer_0[1423] & layer_0[1126]); 
    assign out[1727] = layer_0[249] ^ layer_0[697]; 
    assign out[1728] = ~layer_0[90]; 
    assign out[1729] = layer_0[1135]; 
    assign out[1730] = layer_0[864] & ~layer_0[1065]; 
    assign out[1731] = layer_0[2253] | layer_0[2193]; 
    assign out[1732] = layer_0[786]; 
    assign out[1733] = layer_0[1984] & ~layer_0[2373]; 
    assign out[1734] = ~(layer_0[1238] ^ layer_0[2393]); 
    assign out[1735] = ~(layer_0[1027] ^ layer_0[826]); 
    assign out[1736] = ~(layer_0[193] ^ layer_0[1582]); 
    assign out[1737] = ~layer_0[653]; 
    assign out[1738] = layer_0[921] & ~layer_0[2541]; 
    assign out[1739] = layer_0[2144] | layer_0[339]; 
    assign out[1740] = layer_0[2549] & ~layer_0[1562]; 
    assign out[1741] = layer_0[1984]; 
    assign out[1742] = ~layer_0[914] | (layer_0[914] & layer_0[1692]); 
    assign out[1743] = ~layer_0[512]; 
    assign out[1744] = ~(layer_0[1422] | layer_0[1501]); 
    assign out[1745] = ~layer_0[1260]; 
    assign out[1746] = ~layer_0[1273]; 
    assign out[1747] = layer_0[2148] & layer_0[2018]; 
    assign out[1748] = layer_0[2171] ^ layer_0[2114]; 
    assign out[1749] = ~layer_0[310]; 
    assign out[1750] = ~(layer_0[2342] ^ layer_0[54]); 
    assign out[1751] = ~(layer_0[992] ^ layer_0[795]); 
    assign out[1752] = layer_0[2173]; 
    assign out[1753] = layer_0[1330] & ~layer_0[1972]; 
    assign out[1754] = ~layer_0[2350]; 
    assign out[1755] = ~layer_0[2292] | (layer_0[2292] & layer_0[615]); 
    assign out[1756] = layer_0[2284] ^ layer_0[1596]; 
    assign out[1757] = layer_0[177]; 
    assign out[1758] = layer_0[392] ^ layer_0[1266]; 
    assign out[1759] = layer_0[572]; 
    assign out[1760] = layer_0[2526] ^ layer_0[947]; 
    assign out[1761] = layer_0[119]; 
    assign out[1762] = ~layer_0[1762]; 
    assign out[1763] = ~layer_0[1349]; 
    assign out[1764] = ~layer_0[713]; 
    assign out[1765] = ~layer_0[701]; 
    assign out[1766] = layer_0[1979] ^ layer_0[518]; 
    assign out[1767] = ~(layer_0[622] | layer_0[1751]); 
    assign out[1768] = ~layer_0[2142] | (layer_0[2253] & layer_0[2142]); 
    assign out[1769] = ~layer_0[1970]; 
    assign out[1770] = ~(layer_0[1001] | layer_0[1796]); 
    assign out[1771] = layer_0[438] & layer_0[5]; 
    assign out[1772] = layer_0[1496] & ~layer_0[173]; 
    assign out[1773] = ~layer_0[917]; 
    assign out[1774] = layer_0[2340]; 
    assign out[1775] = ~layer_0[522] | (layer_0[522] & layer_0[800]); 
    assign out[1776] = ~(layer_0[1484] | layer_0[193]); 
    assign out[1777] = layer_0[1097] & ~layer_0[101]; 
    assign out[1778] = layer_0[618] & ~layer_0[2453]; 
    assign out[1779] = layer_0[1139]; 
    assign out[1780] = layer_0[503] ^ layer_0[2468]; 
    assign out[1781] = layer_0[1607]; 
    assign out[1782] = layer_0[2437] & layer_0[1804]; 
    assign out[1783] = layer_0[343] ^ layer_0[904]; 
    assign out[1784] = layer_0[221] & layer_0[384]; 
    assign out[1785] = layer_0[2161] & layer_0[219]; 
    assign out[1786] = layer_0[462] & ~layer_0[2341]; 
    assign out[1787] = layer_0[1929] ^ layer_0[847]; 
    assign out[1788] = layer_0[2528] & ~layer_0[1609]; 
    assign out[1789] = layer_0[2161] & ~layer_0[732]; 
    assign out[1790] = ~layer_0[1731]; 
    assign out[1791] = layer_0[1533] & ~layer_0[2554]; 
    assign out[1792] = layer_0[70]; 
    assign out[1793] = ~(layer_0[1952] | layer_0[218]); 
    assign out[1794] = ~(layer_0[1727] ^ layer_0[965]); 
    assign out[1795] = ~layer_0[763]; 
    assign out[1796] = layer_0[910] & ~layer_0[1289]; 
    assign out[1797] = layer_0[205]; 
    assign out[1798] = ~(layer_0[542] | layer_0[2374]); 
    assign out[1799] = layer_0[1896] & layer_0[2314]; 
    assign out[1800] = layer_0[914] | layer_0[256]; 
    assign out[1801] = layer_0[645] ^ layer_0[1567]; 
    assign out[1802] = ~layer_0[443]; 
    assign out[1803] = ~layer_0[496] | (layer_0[496] & layer_0[638]); 
    assign out[1804] = ~(layer_0[822] & layer_0[2109]); 
    assign out[1805] = layer_0[1257] ^ layer_0[1520]; 
    assign out[1806] = layer_0[2085]; 
    assign out[1807] = layer_0[1818]; 
    assign out[1808] = ~layer_0[1308]; 
    assign out[1809] = layer_0[1608] & layer_0[2404]; 
    assign out[1810] = layer_0[1950] ^ layer_0[1942]; 
    assign out[1811] = layer_0[636]; 
    assign out[1812] = layer_0[2127] & ~layer_0[763]; 
    assign out[1813] = layer_0[2223] & ~layer_0[2256]; 
    assign out[1814] = layer_0[2318] | layer_0[111]; 
    assign out[1815] = layer_0[1921]; 
    assign out[1816] = layer_0[2007] & ~layer_0[1345]; 
    assign out[1817] = layer_0[2431]; 
    assign out[1818] = layer_0[1785] & ~layer_0[1483]; 
    assign out[1819] = layer_0[1998]; 
    assign out[1820] = layer_0[1186] & layer_0[1341]; 
    assign out[1821] = ~layer_0[1854]; 
    assign out[1822] = ~(layer_0[259] ^ layer_0[2094]); 
    assign out[1823] = layer_0[1862] ^ layer_0[2286]; 
    assign out[1824] = layer_0[1785] & ~layer_0[1824]; 
    assign out[1825] = ~(layer_0[2166] | layer_0[75]); 
    assign out[1826] = ~layer_0[1323]; 
    assign out[1827] = ~layer_0[1330]; 
    assign out[1828] = layer_0[40]; 
    assign out[1829] = layer_0[1702] ^ layer_0[2243]; 
    assign out[1830] = ~layer_0[482]; 
    assign out[1831] = layer_0[655] ^ layer_0[2124]; 
    assign out[1832] = ~layer_0[1618] | (layer_0[1618] & layer_0[1051]); 
    assign out[1833] = layer_0[1764] & ~layer_0[2309]; 
    assign out[1834] = ~(layer_0[1060] | layer_0[1781]); 
    assign out[1835] = layer_0[2403] ^ layer_0[808]; 
    assign out[1836] = layer_0[1210] & ~layer_0[1031]; 
    assign out[1837] = ~layer_0[1042]; 
    assign out[1838] = ~layer_0[2467]; 
    assign out[1839] = layer_0[2276]; 
    assign out[1840] = layer_0[282] & ~layer_0[639]; 
    assign out[1841] = ~(layer_0[2171] ^ layer_0[2543]); 
    assign out[1842] = ~(layer_0[260] ^ layer_0[631]); 
    assign out[1843] = layer_0[90] & ~layer_0[357]; 
    assign out[1844] = layer_0[826] | layer_0[365]; 
    assign out[1845] = layer_0[964] & layer_0[675]; 
    assign out[1846] = layer_0[456] & layer_0[2016]; 
    assign out[1847] = layer_0[2453]; 
    assign out[1848] = ~(layer_0[2018] | layer_0[164]); 
    assign out[1849] = ~layer_0[1883]; 
    assign out[1850] = ~(layer_0[610] | layer_0[781]); 
    assign out[1851] = layer_0[94] & ~layer_0[1604]; 
    assign out[1852] = layer_0[1100] & ~layer_0[1825]; 
    assign out[1853] = ~layer_0[539] | (layer_0[539] & layer_0[2276]); 
    assign out[1854] = ~layer_0[2294] | (layer_0[2294] & layer_0[2384]); 
    assign out[1855] = ~(layer_0[2076] | layer_0[2441]); 
    assign out[1856] = layer_0[1830] ^ layer_0[2062]; 
    assign out[1857] = layer_0[383] & ~layer_0[1238]; 
    assign out[1858] = layer_0[814]; 
    assign out[1859] = layer_0[2157]; 
    assign out[1860] = layer_0[651] | layer_0[1104]; 
    assign out[1861] = layer_0[2122] ^ layer_0[1342]; 
    assign out[1862] = ~layer_0[376]; 
    assign out[1863] = ~layer_0[307]; 
    assign out[1864] = layer_0[1753]; 
    assign out[1865] = layer_0[1720]; 
    assign out[1866] = ~layer_0[1854]; 
    assign out[1867] = layer_0[1941]; 
    assign out[1868] = layer_0[2484]; 
    assign out[1869] = layer_0[1931] & ~layer_0[1225]; 
    assign out[1870] = ~layer_0[218] | (layer_0[634] & layer_0[218]); 
    assign out[1871] = layer_0[2258] ^ layer_0[1391]; 
    assign out[1872] = ~layer_0[2072]; 
    assign out[1873] = ~(layer_0[2479] ^ layer_0[1686]); 
    assign out[1874] = layer_0[1828] | layer_0[2536]; 
    assign out[1875] = ~(layer_0[2102] ^ layer_0[1380]); 
    assign out[1876] = ~(layer_0[1471] ^ layer_0[849]); 
    assign out[1877] = ~layer_0[921]; 
    assign out[1878] = layer_0[1679] & layer_0[1177]; 
    assign out[1879] = layer_0[226] & ~layer_0[1083]; 
    assign out[1880] = layer_0[2056]; 
    assign out[1881] = layer_0[796]; 
    assign out[1882] = layer_0[862]; 
    assign out[1883] = layer_0[901] & layer_0[1720]; 
    assign out[1884] = ~layer_0[537]; 
    assign out[1885] = ~(layer_0[708] | layer_0[1841]); 
    assign out[1886] = layer_0[1821] ^ layer_0[697]; 
    assign out[1887] = ~layer_0[2027] | (layer_0[2027] & layer_0[675]); 
    assign out[1888] = layer_0[2211]; 
    assign out[1889] = layer_0[2337] ^ layer_0[2325]; 
    assign out[1890] = ~(layer_0[1426] ^ layer_0[1125]); 
    assign out[1891] = ~(layer_0[1469] ^ layer_0[2265]); 
    assign out[1892] = ~layer_0[1584] | (layer_0[957] & layer_0[1584]); 
    assign out[1893] = ~(layer_0[2467] | layer_0[857]); 
    assign out[1894] = ~(layer_0[2197] ^ layer_0[2289]); 
    assign out[1895] = ~(layer_0[1647] | layer_0[1225]); 
    assign out[1896] = ~layer_0[825]; 
    assign out[1897] = ~layer_0[5]; 
    assign out[1898] = layer_0[592]; 
    assign out[1899] = ~(layer_0[501] ^ layer_0[1670]); 
    assign out[1900] = ~layer_0[921]; 
    assign out[1901] = layer_0[1635] & layer_0[461]; 
    assign out[1902] = ~layer_0[2089]; 
    assign out[1903] = ~layer_0[848] | (layer_0[388] & layer_0[848]); 
    assign out[1904] = ~layer_0[359]; 
    assign out[1905] = ~(layer_0[1854] | layer_0[1369]); 
    assign out[1906] = ~layer_0[700]; 
    assign out[1907] = ~(layer_0[1456] | layer_0[386]); 
    assign out[1908] = layer_0[1141] & layer_0[2154]; 
    assign out[1909] = layer_0[508]; 
    assign out[1910] = layer_0[1493] & ~layer_0[2053]; 
    assign out[1911] = ~(layer_0[1867] | layer_0[1369]); 
    assign out[1912] = layer_0[558] & ~layer_0[1356]; 
    assign out[1913] = layer_0[108] & layer_0[239]; 
    assign out[1914] = layer_0[2246] ^ layer_0[2477]; 
    assign out[1915] = layer_0[145] & ~layer_0[425]; 
    assign out[1916] = layer_0[1015] & ~layer_0[9]; 
    assign out[1917] = ~layer_0[1847]; 
    assign out[1918] = ~(layer_0[207] | layer_0[478]); 
    assign out[1919] = layer_0[842] & ~layer_0[1867]; 
    assign out[1920] = ~(layer_0[2274] ^ layer_0[2170]); 
    assign out[1921] = layer_0[1325] | layer_0[990]; 
    assign out[1922] = ~(layer_0[590] ^ layer_0[1083]); 
    assign out[1923] = ~layer_0[2003]; 
    assign out[1924] = layer_0[1673] ^ layer_0[2080]; 
    assign out[1925] = layer_0[1709] & layer_0[1231]; 
    assign out[1926] = layer_0[847] ^ layer_0[1088]; 
    assign out[1927] = layer_0[1347]; 
    assign out[1928] = ~(layer_0[1244] ^ layer_0[905]); 
    assign out[1929] = layer_0[939]; 
    assign out[1930] = layer_0[48] & layer_0[2211]; 
    assign out[1931] = ~layer_0[1850]; 
    assign out[1932] = ~layer_0[1924]; 
    assign out[1933] = ~(layer_0[398] ^ layer_0[1102]); 
    assign out[1934] = layer_0[1944] ^ layer_0[2042]; 
    assign out[1935] = layer_0[1241] & layer_0[107]; 
    assign out[1936] = layer_0[2314]; 
    assign out[1937] = layer_0[2496] & ~layer_0[2144]; 
    assign out[1938] = layer_0[927] ^ layer_0[2471]; 
    assign out[1939] = ~layer_0[496]; 
    assign out[1940] = layer_0[1015] & layer_0[1347]; 
    assign out[1941] = ~(layer_0[1193] ^ layer_0[1686]); 
    assign out[1942] = layer_0[1492] & ~layer_0[2285]; 
    assign out[1943] = ~(layer_0[2365] ^ layer_0[2009]); 
    assign out[1944] = layer_0[2157]; 
    assign out[1945] = layer_0[1618] ^ layer_0[144]; 
    assign out[1946] = layer_0[1164]; 
    assign out[1947] = layer_0[2498] ^ layer_0[1718]; 
    assign out[1948] = layer_0[934] & layer_0[2367]; 
    assign out[1949] = layer_0[671]; 
    assign out[1950] = ~(layer_0[568] ^ layer_0[1526]); 
    assign out[1951] = ~layer_0[1195] | (layer_0[1195] & layer_0[983]); 
    assign out[1952] = layer_0[346] & ~layer_0[1757]; 
    assign out[1953] = layer_0[1445] & ~layer_0[2497]; 
    assign out[1954] = layer_0[1869] & ~layer_0[840]; 
    assign out[1955] = ~layer_0[1326]; 
    assign out[1956] = layer_0[389] ^ layer_0[2329]; 
    assign out[1957] = layer_0[2476] & layer_0[388]; 
    assign out[1958] = ~(layer_0[1085] ^ layer_0[672]); 
    assign out[1959] = ~(layer_0[1134] | layer_0[372]); 
    assign out[1960] = layer_0[741]; 
    assign out[1961] = ~(layer_0[1403] ^ layer_0[562]); 
    assign out[1962] = layer_0[606] | layer_0[26]; 
    assign out[1963] = ~layer_0[926] | (layer_0[926] & layer_0[903]); 
    assign out[1964] = ~layer_0[2353]; 
    assign out[1965] = ~layer_0[1331]; 
    assign out[1966] = layer_0[1720] ^ layer_0[1129]; 
    assign out[1967] = layer_0[1921] & ~layer_0[478]; 
    assign out[1968] = layer_0[1408] ^ layer_0[1979]; 
    assign out[1969] = ~layer_0[1193] | (layer_0[1608] & layer_0[1193]); 
    assign out[1970] = layer_0[2381] & ~layer_0[2386]; 
    assign out[1971] = layer_0[616] & ~layer_0[955]; 
    assign out[1972] = ~(layer_0[1583] & layer_0[1666]); 
    assign out[1973] = layer_0[930] & ~layer_0[496]; 
    assign out[1974] = ~(layer_0[138] ^ layer_0[405]); 
    assign out[1975] = ~(layer_0[821] ^ layer_0[1683]); 
    assign out[1976] = layer_0[727] ^ layer_0[884]; 
    assign out[1977] = ~layer_0[1378]; 
    assign out[1978] = layer_0[1572] & ~layer_0[2317]; 
    assign out[1979] = ~(layer_0[1669] | layer_0[2072]); 
    assign out[1980] = ~layer_0[1587]; 
    assign out[1981] = ~layer_0[2374]; 
    assign out[1982] = ~(layer_0[1458] | layer_0[551]); 
    assign out[1983] = layer_0[321]; 
    assign out[1984] = layer_0[1700] & ~layer_0[438]; 
    assign out[1985] = layer_0[533] ^ layer_0[2415]; 
    assign out[1986] = layer_0[25]; 
    assign out[1987] = layer_0[1176] & ~layer_0[1731]; 
    assign out[1988] = ~layer_0[1886]; 
    assign out[1989] = layer_0[528] ^ layer_0[232]; 
    assign out[1990] = ~layer_0[140]; 
    assign out[1991] = ~layer_0[496]; 
    assign out[1992] = layer_0[2512]; 
    assign out[1993] = ~layer_0[2374]; 
    assign out[1994] = layer_0[1772] ^ layer_0[1510]; 
    assign out[1995] = layer_0[346]; 
    assign out[1996] = ~(layer_0[722] ^ layer_0[1125]); 
    assign out[1997] = ~(layer_0[2113] | layer_0[386]); 
    assign out[1998] = layer_0[1121] ^ layer_0[1339]; 
    assign out[1999] = ~(layer_0[2028] | layer_0[1461]); 
    assign out[2000] = layer_0[1323] ^ layer_0[1244]; 
    assign out[2001] = layer_0[787] & ~layer_0[427]; 
    assign out[2002] = ~layer_0[143]; 
    assign out[2003] = layer_0[2016] & ~layer_0[1323]; 
    assign out[2004] = layer_0[391]; 
    assign out[2005] = ~(layer_0[1680] | layer_0[1554]); 
    assign out[2006] = layer_0[637] & ~layer_0[443]; 
    assign out[2007] = layer_0[396] & layer_0[882]; 
    assign out[2008] = layer_0[1469]; 
    assign out[2009] = layer_0[254] ^ layer_0[1104]; 
    assign out[2010] = layer_0[1695]; 
    assign out[2011] = ~(layer_0[496] | layer_0[2018]); 
    assign out[2012] = layer_0[1059] & layer_0[2161]; 
    assign out[2013] = ~layer_0[1103] | (layer_0[1902] & layer_0[1103]); 
    assign out[2014] = layer_0[2134] ^ layer_0[344]; 
    assign out[2015] = ~(layer_0[2273] ^ layer_0[1554]); 
    assign out[2016] = layer_0[145]; 
    assign out[2017] = ~layer_0[1847]; 
    assign out[2018] = ~layer_0[1034]; 
    assign out[2019] = ~(layer_0[1118] & layer_0[1583]); 
    assign out[2020] = layer_0[2205] ^ layer_0[101]; 
    assign out[2021] = layer_0[1625]; 
    assign out[2022] = ~(layer_0[218] & layer_0[2012]); 
    assign out[2023] = layer_0[1463] & ~layer_0[2557]; 
    assign out[2024] = ~(layer_0[117] ^ layer_0[483]); 
    assign out[2025] = layer_0[77] ^ layer_0[1933]; 
    assign out[2026] = ~(layer_0[1841] ^ layer_0[2160]); 
    assign out[2027] = ~layer_0[866]; 
    assign out[2028] = layer_0[205]; 
    assign out[2029] = layer_0[709] | layer_0[914]; 
    assign out[2030] = layer_0[1553] & layer_0[2367]; 
    assign out[2031] = ~(layer_0[1880] ^ layer_0[728]); 
    assign out[2032] = ~(layer_0[1443] ^ layer_0[1417]); 
    assign out[2033] = ~layer_0[2132] | (layer_0[2132] & layer_0[198]); 
    assign out[2034] = ~(layer_0[532] ^ layer_0[1578]); 
    assign out[2035] = ~(layer_0[2342] ^ layer_0[2336]); 
    assign out[2036] = layer_0[2225]; 
    assign out[2037] = layer_0[2126] | layer_0[2181]; 
    assign out[2038] = layer_0[91] ^ layer_0[1368]; 
    assign out[2039] = ~layer_0[1321] | (layer_0[2543] & layer_0[1321]); 
    assign out[2040] = ~(layer_0[1476] ^ layer_0[2068]); 
    assign out[2041] = layer_0[739]; 
    assign out[2042] = ~(layer_0[1626] ^ layer_0[2034]); 
    assign out[2043] = layer_0[1845]; 
    assign out[2044] = ~layer_0[117]; 
    assign out[2045] = ~(layer_0[2088] ^ layer_0[2043]); 
    assign out[2046] = ~layer_0[1356]; 
    assign out[2047] = layer_0[568] ^ layer_0[472]; 
    assign out[2048] = ~layer_0[1048]; 
    assign out[2049] = layer_0[714]; 
    assign out[2050] = ~layer_0[2527]; 
    assign out[2051] = ~(layer_0[404] ^ layer_0[1520]); 
    assign out[2052] = layer_0[1563] & layer_0[1952]; 
    assign out[2053] = layer_0[1934]; 
    assign out[2054] = layer_0[737] | layer_0[2345]; 
    assign out[2055] = ~(layer_0[2472] ^ layer_0[2314]); 
    assign out[2056] = ~(layer_0[1463] ^ layer_0[1191]); 
    assign out[2057] = layer_0[159] & ~layer_0[960]; 
    assign out[2058] = layer_0[568] ^ layer_0[2501]; 
    assign out[2059] = layer_0[1248] | layer_0[887]; 
    assign out[2060] = layer_0[233] ^ layer_0[1707]; 
    assign out[2061] = layer_0[580] | layer_0[159]; 
    assign out[2062] = ~(layer_0[1950] ^ layer_0[2124]); 
    assign out[2063] = layer_0[1204] ^ layer_0[1879]; 
    assign out[2064] = layer_0[2535] & ~layer_0[1480]; 
    assign out[2065] = ~layer_0[860] | (layer_0[1862] & layer_0[860]); 
    assign out[2066] = layer_0[1522] ^ layer_0[2341]; 
    assign out[2067] = ~(layer_0[529] ^ layer_0[846]); 
    assign out[2068] = layer_0[2226] ^ layer_0[725]; 
    assign out[2069] = layer_0[688]; 
    assign out[2070] = ~(layer_0[341] ^ layer_0[728]); 
    assign out[2071] = layer_0[1881] & ~layer_0[104]; 
    assign out[2072] = layer_0[1673]; 
    assign out[2073] = ~layer_0[752]; 
    assign out[2074] = layer_0[589] & layer_0[1708]; 
    assign out[2075] = ~(layer_0[864] | layer_0[393]); 
    assign out[2076] = layer_0[340] & ~layer_0[541]; 
    assign out[2077] = ~layer_0[999]; 
    assign out[2078] = ~(layer_0[1661] ^ layer_0[1734]); 
    assign out[2079] = layer_0[1491] & ~layer_0[232]; 
    assign out[2080] = ~layer_0[449]; 
    assign out[2081] = layer_0[2206]; 
    assign out[2082] = ~(layer_0[389] ^ layer_0[1134]); 
    assign out[2083] = ~layer_0[1769]; 
    assign out[2084] = ~(layer_0[1187] ^ layer_0[2369]); 
    assign out[2085] = layer_0[1435]; 
    assign out[2086] = layer_0[1678] ^ layer_0[2425]; 
    assign out[2087] = ~layer_0[56]; 
    assign out[2088] = ~(layer_0[939] | layer_0[1115]); 
    assign out[2089] = layer_0[1506]; 
    assign out[2090] = ~(layer_0[1327] ^ layer_0[687]); 
    assign out[2091] = ~(layer_0[576] ^ layer_0[1076]); 
    assign out[2092] = ~(layer_0[2094] ^ layer_0[985]); 
    assign out[2093] = layer_0[1956]; 
    assign out[2094] = ~(layer_0[724] ^ layer_0[798]); 
    assign out[2095] = ~layer_0[2250]; 
    assign out[2096] = layer_0[2347] ^ layer_0[1128]; 
    assign out[2097] = ~layer_0[2176]; 
    assign out[2098] = layer_0[1083] & ~layer_0[1973]; 
    assign out[2099] = layer_0[589] | layer_0[519]; 
    assign out[2100] = layer_0[974] & ~layer_0[993]; 
    assign out[2101] = ~(layer_0[623] ^ layer_0[1016]); 
    assign out[2102] = layer_0[2301]; 
    assign out[2103] = ~layer_0[1973] | (layer_0[2094] & layer_0[1973]); 
    assign out[2104] = layer_0[2076] ^ layer_0[1758]; 
    assign out[2105] = ~layer_0[2042] | (layer_0[1258] & layer_0[2042]); 
    assign out[2106] = layer_0[1402] ^ layer_0[1713]; 
    assign out[2107] = layer_0[1258]; 
    assign out[2108] = ~layer_0[2445]; 
    assign out[2109] = layer_0[1447] & ~layer_0[449]; 
    assign out[2110] = layer_0[1311]; 
    assign out[2111] = ~(layer_0[2040] ^ layer_0[2546]); 
    assign out[2112] = ~layer_0[2491]; 
    assign out[2113] = layer_0[2107]; 
    assign out[2114] = ~(layer_0[1424] ^ layer_0[1131]); 
    assign out[2115] = ~(layer_0[2305] & layer_0[889]); 
    assign out[2116] = ~(layer_0[662] ^ layer_0[122]); 
    assign out[2117] = layer_0[1799]; 
    assign out[2118] = ~(layer_0[1498] ^ layer_0[993]); 
    assign out[2119] = ~layer_0[1482]; 
    assign out[2120] = ~layer_0[788] | (layer_0[1524] & layer_0[788]); 
    assign out[2121] = layer_0[422] ^ layer_0[720]; 
    assign out[2122] = ~(layer_0[1630] & layer_0[1693]); 
    assign out[2123] = layer_0[351] ^ layer_0[468]; 
    assign out[2124] = ~(layer_0[2154] ^ layer_0[1143]); 
    assign out[2125] = ~layer_0[1480] | (layer_0[1847] & layer_0[1480]); 
    assign out[2126] = ~(layer_0[232] & layer_0[1795]); 
    assign out[2127] = layer_0[239] ^ layer_0[1269]; 
    assign out[2128] = ~(layer_0[1978] ^ layer_0[423]); 
    assign out[2129] = layer_0[809] ^ layer_0[1454]; 
    assign out[2130] = ~layer_0[2421] | (layer_0[2421] & layer_0[151]); 
    assign out[2131] = ~(layer_0[2337] & layer_0[962]); 
    assign out[2132] = layer_0[2235]; 
    assign out[2133] = ~layer_0[1618] | (layer_0[1618] & layer_0[1317]); 
    assign out[2134] = layer_0[19] ^ layer_0[973]; 
    assign out[2135] = ~(layer_0[1973] & layer_0[352]); 
    assign out[2136] = layer_0[406]; 
    assign out[2137] = layer_0[2500] | layer_0[1858]; 
    assign out[2138] = ~layer_0[1482]; 
    assign out[2139] = layer_0[534]; 
    assign out[2140] = layer_0[1057] ^ layer_0[873]; 
    assign out[2141] = ~layer_0[647] | (layer_0[647] & layer_0[1744]); 
    assign out[2142] = layer_0[454] ^ layer_0[1419]; 
    assign out[2143] = layer_0[1525]; 
    assign out[2144] = layer_0[944] ^ layer_0[1698]; 
    assign out[2145] = layer_0[1401] & ~layer_0[75]; 
    assign out[2146] = ~layer_0[741]; 
    assign out[2147] = ~layer_0[1380]; 
    assign out[2148] = ~(layer_0[1594] & layer_0[2332]); 
    assign out[2149] = layer_0[2468] & ~layer_0[2499]; 
    assign out[2150] = layer_0[1986]; 
    assign out[2151] = layer_0[1216]; 
    assign out[2152] = layer_0[1422]; 
    assign out[2153] = ~layer_0[37] | (layer_0[340] & layer_0[37]); 
    assign out[2154] = layer_0[546] ^ layer_0[972]; 
    assign out[2155] = ~(layer_0[2505] ^ layer_0[1246]); 
    assign out[2156] = layer_0[2258] & ~layer_0[2336]; 
    assign out[2157] = layer_0[896] & layer_0[594]; 
    assign out[2158] = ~(layer_0[702] ^ layer_0[792]); 
    assign out[2159] = ~layer_0[720]; 
    assign out[2160] = layer_0[1726]; 
    assign out[2161] = ~layer_0[592]; 
    assign out[2162] = ~layer_0[2238]; 
    assign out[2163] = layer_0[496] & ~layer_0[1865]; 
    assign out[2164] = ~layer_0[1098]; 
    assign out[2165] = ~(layer_0[78] ^ layer_0[1943]); 
    assign out[2166] = layer_0[473] ^ layer_0[1970]; 
    assign out[2167] = ~(layer_0[51] | layer_0[572]); 
    assign out[2168] = layer_0[1626] & ~layer_0[769]; 
    assign out[2169] = ~layer_0[2091]; 
    assign out[2170] = layer_0[364] ^ layer_0[2021]; 
    assign out[2171] = ~(layer_0[810] ^ layer_0[861]); 
    assign out[2172] = ~(layer_0[1451] ^ layer_0[550]); 
    assign out[2173] = ~(layer_0[371] ^ layer_0[605]); 
    assign out[2174] = ~(layer_0[1385] ^ layer_0[823]); 
    assign out[2175] = ~layer_0[1540]; 
    assign out[2176] = layer_0[1736]; 
    assign out[2177] = layer_0[1448]; 
    assign out[2178] = ~(layer_0[885] ^ layer_0[1842]); 
    assign out[2179] = ~(layer_0[890] & layer_0[249]); 
    assign out[2180] = ~layer_0[636] | (layer_0[274] & layer_0[636]); 
    assign out[2181] = layer_0[1483] & ~layer_0[2312]; 
    assign out[2182] = ~(layer_0[389] | layer_0[1429]); 
    assign out[2183] = ~(layer_0[634] ^ layer_0[970]); 
    assign out[2184] = layer_0[781] ^ layer_0[373]; 
    assign out[2185] = ~(layer_0[516] | layer_0[908]); 
    assign out[2186] = ~(layer_0[2202] ^ layer_0[2246]); 
    assign out[2187] = ~(layer_0[1235] ^ layer_0[850]); 
    assign out[2188] = layer_0[1914] & ~layer_0[1440]; 
    assign out[2189] = ~(layer_0[852] | layer_0[997]); 
    assign out[2190] = ~layer_0[1923]; 
    assign out[2191] = ~(layer_0[2526] ^ layer_0[1471]); 
    assign out[2192] = ~(layer_0[1897] ^ layer_0[147]); 
    assign out[2193] = ~layer_0[1617]; 
    assign out[2194] = ~layer_0[97]; 
    assign out[2195] = layer_0[1574] ^ layer_0[2057]; 
    assign out[2196] = layer_0[2049]; 
    assign out[2197] = layer_0[1414] ^ layer_0[1718]; 
    assign out[2198] = layer_0[1522] ^ layer_0[298]; 
    assign out[2199] = ~(layer_0[1410] ^ layer_0[2306]); 
    assign out[2200] = ~(layer_0[2297] ^ layer_0[1016]); 
    assign out[2201] = layer_0[395] ^ layer_0[2399]; 
    assign out[2202] = ~(layer_0[84] ^ layer_0[341]); 
    assign out[2203] = layer_0[2326] ^ layer_0[592]; 
    assign out[2204] = ~(layer_0[804] | layer_0[380]); 
    assign out[2205] = layer_0[1934] & ~layer_0[1945]; 
    assign out[2206] = layer_0[688]; 
    assign out[2207] = layer_0[1462] & layer_0[816]; 
    assign out[2208] = layer_0[696]; 
    assign out[2209] = ~layer_0[417] | (layer_0[1452] & layer_0[417]); 
    assign out[2210] = ~layer_0[1097]; 
    assign out[2211] = ~(layer_0[2089] ^ layer_0[68]); 
    assign out[2212] = layer_0[2012] ^ layer_0[727]; 
    assign out[2213] = ~layer_0[1613] | (layer_0[1613] & layer_0[519]); 
    assign out[2214] = ~(layer_0[395] ^ layer_0[2096]); 
    assign out[2215] = layer_0[2362] ^ layer_0[1003]; 
    assign out[2216] = ~(layer_0[1987] ^ layer_0[1287]); 
    assign out[2217] = layer_0[231] ^ layer_0[2419]; 
    assign out[2218] = ~layer_0[1534] | (layer_0[1534] & layer_0[2535]); 
    assign out[2219] = layer_0[1799]; 
    assign out[2220] = layer_0[537] & ~layer_0[962]; 
    assign out[2221] = ~(layer_0[507] ^ layer_0[751]); 
    assign out[2222] = ~layer_0[1594] | (layer_0[1855] & layer_0[1594]); 
    assign out[2223] = layer_0[521] ^ layer_0[678]; 
    assign out[2224] = layer_0[735] ^ layer_0[1909]; 
    assign out[2225] = layer_0[901]; 
    assign out[2226] = ~layer_0[1683]; 
    assign out[2227] = layer_0[714]; 
    assign out[2228] = ~layer_0[2035]; 
    assign out[2229] = ~layer_0[1091]; 
    assign out[2230] = layer_0[1024] ^ layer_0[1824]; 
    assign out[2231] = layer_0[2558]; 
    assign out[2232] = ~layer_0[790]; 
    assign out[2233] = layer_0[717]; 
    assign out[2234] = ~layer_0[385] | (layer_0[823] & layer_0[385]); 
    assign out[2235] = ~layer_0[644]; 
    assign out[2236] = layer_0[2193] ^ layer_0[2108]; 
    assign out[2237] = layer_0[263] ^ layer_0[21]; 
    assign out[2238] = ~(layer_0[1055] ^ layer_0[477]); 
    assign out[2239] = layer_0[451] | layer_0[492]; 
    assign out[2240] = layer_0[2095] | layer_0[2535]; 
    assign out[2241] = ~layer_0[2143]; 
    assign out[2242] = ~(layer_0[845] & layer_0[17]); 
    assign out[2243] = ~(layer_0[2233] ^ layer_0[2531]); 
    assign out[2244] = layer_0[1379] & layer_0[133]; 
    assign out[2245] = layer_0[1242]; 
    assign out[2246] = layer_0[1799]; 
    assign out[2247] = ~(layer_0[2022] | layer_0[2318]); 
    assign out[2248] = layer_0[1038] | layer_0[1275]; 
    assign out[2249] = ~(layer_0[1700] ^ layer_0[163]); 
    assign out[2250] = layer_0[1845]; 
    assign out[2251] = layer_0[1708] | layer_0[1298]; 
    assign out[2252] = layer_0[2380] ^ layer_0[1649]; 
    assign out[2253] = ~(layer_0[2245] ^ layer_0[692]); 
    assign out[2254] = ~(layer_0[2462] ^ layer_0[2154]); 
    assign out[2255] = layer_0[2234] ^ layer_0[671]; 
    assign out[2256] = ~layer_0[1423]; 
    assign out[2257] = ~layer_0[2318]; 
    assign out[2258] = ~layer_0[1514]; 
    assign out[2259] = ~(layer_0[576] ^ layer_0[1712]); 
    assign out[2260] = ~layer_0[1377] | (layer_0[1377] & layer_0[216]); 
    assign out[2261] = layer_0[1379] & ~layer_0[1617]; 
    assign out[2262] = ~(layer_0[324] ^ layer_0[1350]); 
    assign out[2263] = layer_0[1196] & ~layer_0[543]; 
    assign out[2264] = ~(layer_0[13] ^ layer_0[699]); 
    assign out[2265] = layer_0[1598] | layer_0[1506]; 
    assign out[2266] = layer_0[971] ^ layer_0[947]; 
    assign out[2267] = ~(layer_0[1624] ^ layer_0[1160]); 
    assign out[2268] = layer_0[1173]; 
    assign out[2269] = ~layer_0[249]; 
    assign out[2270] = ~(layer_0[433] ^ layer_0[1644]); 
    assign out[2271] = layer_0[2141] ^ layer_0[2094]; 
    assign out[2272] = ~layer_0[2358] | (layer_0[1375] & layer_0[2358]); 
    assign out[2273] = ~(layer_0[2528] ^ layer_0[1240]); 
    assign out[2274] = ~(layer_0[1594] & layer_0[463]); 
    assign out[2275] = ~(layer_0[360] ^ layer_0[892]); 
    assign out[2276] = ~layer_0[1987] | (layer_0[1987] & layer_0[2415]); 
    assign out[2277] = ~(layer_0[2553] ^ layer_0[28]); 
    assign out[2278] = layer_0[1289]; 
    assign out[2279] = layer_0[2002] | layer_0[2354]; 
    assign out[2280] = ~(layer_0[37] | layer_0[1221]); 
    assign out[2281] = layer_0[171] ^ layer_0[164]; 
    assign out[2282] = layer_0[59] ^ layer_0[2416]; 
    assign out[2283] = layer_0[63]; 
    assign out[2284] = layer_0[1919] ^ layer_0[1815]; 
    assign out[2285] = ~layer_0[1640] | (layer_0[715] & layer_0[1640]); 
    assign out[2286] = layer_0[406]; 
    assign out[2287] = layer_0[1019] ^ layer_0[648]; 
    assign out[2288] = layer_0[1462] | layer_0[1438]; 
    assign out[2289] = layer_0[1422]; 
    assign out[2290] = layer_0[2212] ^ layer_0[1791]; 
    assign out[2291] = ~(layer_0[701] ^ layer_0[1902]); 
    assign out[2292] = ~(layer_0[2233] & layer_0[1205]); 
    assign out[2293] = ~(layer_0[2112] ^ layer_0[1901]); 
    assign out[2294] = ~layer_0[1720] | (layer_0[1720] & layer_0[2053]); 
    assign out[2295] = layer_0[1611]; 
    assign out[2296] = layer_0[1296]; 
    assign out[2297] = ~layer_0[504]; 
    assign out[2298] = ~(layer_0[1639] | layer_0[1285]); 
    assign out[2299] = layer_0[182] ^ layer_0[1414]; 
    assign out[2300] = ~layer_0[357] | (layer_0[1067] & layer_0[357]); 
    assign out[2301] = layer_0[2178] & layer_0[1622]; 
    assign out[2302] = layer_0[998]; 
    assign out[2303] = layer_0[2413] ^ layer_0[1709]; 
    assign out[2304] = layer_0[2437] | layer_0[289]; 
    assign out[2305] = ~(layer_0[1561] ^ layer_0[807]); 
    assign out[2306] = layer_0[389] & ~layer_0[1515]; 
    assign out[2307] = ~layer_0[1747]; 
    assign out[2308] = ~(layer_0[397] | layer_0[2280]); 
    assign out[2309] = layer_0[847] & ~layer_0[2474]; 
    assign out[2310] = layer_0[1364] ^ layer_0[208]; 
    assign out[2311] = layer_0[868] ^ layer_0[2154]; 
    assign out[2312] = ~layer_0[1588]; 
    assign out[2313] = layer_0[2559] ^ layer_0[276]; 
    assign out[2314] = layer_0[473] & ~layer_0[597]; 
    assign out[2315] = ~layer_0[1327]; 
    assign out[2316] = layer_0[1470] & layer_0[1001]; 
    assign out[2317] = ~layer_0[791]; 
    assign out[2318] = ~(layer_0[343] ^ layer_0[1899]); 
    assign out[2319] = ~(layer_0[2551] | layer_0[555]); 
    assign out[2320] = layer_0[1620] ^ layer_0[1824]; 
    assign out[2321] = layer_0[2322] ^ layer_0[444]; 
    assign out[2322] = ~(layer_0[1941] | layer_0[1365]); 
    assign out[2323] = layer_0[40] ^ layer_0[2247]; 
    assign out[2324] = ~layer_0[160]; 
    assign out[2325] = layer_0[2114] ^ layer_0[688]; 
    assign out[2326] = layer_0[617] ^ layer_0[425]; 
    assign out[2327] = layer_0[2003] & ~layer_0[1193]; 
    assign out[2328] = ~(layer_0[527] ^ layer_0[381]); 
    assign out[2329] = ~(layer_0[697] ^ layer_0[464]); 
    assign out[2330] = layer_0[2156] ^ layer_0[639]; 
    assign out[2331] = ~layer_0[469] | (layer_0[469] & layer_0[2008]); 
    assign out[2332] = layer_0[452] ^ layer_0[1342]; 
    assign out[2333] = ~(layer_0[1437] | layer_0[2239]); 
    assign out[2334] = layer_0[853] & ~layer_0[2214]; 
    assign out[2335] = layer_0[142] & ~layer_0[314]; 
    assign out[2336] = layer_0[1872] ^ layer_0[295]; 
    assign out[2337] = ~(layer_0[610] ^ layer_0[1012]); 
    assign out[2338] = layer_0[821] & layer_0[1165]; 
    assign out[2339] = layer_0[641]; 
    assign out[2340] = ~(layer_0[1309] ^ layer_0[1352]); 
    assign out[2341] = layer_0[998]; 
    assign out[2342] = layer_0[127] & ~layer_0[439]; 
    assign out[2343] = ~(layer_0[1796] | layer_0[845]); 
    assign out[2344] = ~(layer_0[941] | layer_0[1837]); 
    assign out[2345] = ~(layer_0[1340] ^ layer_0[1535]); 
    assign out[2346] = layer_0[1232] & ~layer_0[1799]; 
    assign out[2347] = ~layer_0[431]; 
    assign out[2348] = ~(layer_0[1984] | layer_0[545]); 
    assign out[2349] = ~layer_0[1290] | (layer_0[1290] & layer_0[1546]); 
    assign out[2350] = layer_0[410] & ~layer_0[207]; 
    assign out[2351] = ~(layer_0[1786] | layer_0[772]); 
    assign out[2352] = layer_0[496] ^ layer_0[1544]; 
    assign out[2353] = ~(layer_0[1191] ^ layer_0[50]); 
    assign out[2354] = ~layer_0[1445]; 
    assign out[2355] = ~(layer_0[863] ^ layer_0[334]); 
    assign out[2356] = layer_0[900] & layer_0[1443]; 
    assign out[2357] = layer_0[2338] ^ layer_0[510]; 
    assign out[2358] = layer_0[1970]; 
    assign out[2359] = layer_0[1396] & ~layer_0[535]; 
    assign out[2360] = layer_0[2144]; 
    assign out[2361] = layer_0[2033]; 
    assign out[2362] = layer_0[228] ^ layer_0[1505]; 
    assign out[2363] = layer_0[27] & ~layer_0[586]; 
    assign out[2364] = layer_0[2366] ^ layer_0[2513]; 
    assign out[2365] = layer_0[995] & ~layer_0[1321]; 
    assign out[2366] = layer_0[2206] & ~layer_0[2129]; 
    assign out[2367] = layer_0[2179] & layer_0[532]; 
    assign out[2368] = ~layer_0[674] | (layer_0[2185] & layer_0[674]); 
    assign out[2369] = ~(layer_0[169] ^ layer_0[1498]); 
    assign out[2370] = ~(layer_0[2542] | layer_0[1083]); 
    assign out[2371] = ~(layer_0[2297] | layer_0[1652]); 
    assign out[2372] = layer_0[688] & ~layer_0[50]; 
    assign out[2373] = ~(layer_0[1416] | layer_0[1316]); 
    assign out[2374] = layer_0[2266]; 
    assign out[2375] = ~layer_0[1616]; 
    assign out[2376] = ~(layer_0[673] & layer_0[179]); 
    assign out[2377] = ~layer_0[475]; 
    assign out[2378] = layer_0[300] & ~layer_0[1408]; 
    assign out[2379] = layer_0[2195] ^ layer_0[2027]; 
    assign out[2380] = ~layer_0[211]; 
    assign out[2381] = ~(layer_0[1282] ^ layer_0[952]); 
    assign out[2382] = ~layer_0[2073]; 
    assign out[2383] = layer_0[380]; 
    assign out[2384] = layer_0[2524] ^ layer_0[1666]; 
    assign out[2385] = ~(layer_0[152] ^ layer_0[152]); 
    assign out[2386] = layer_0[793] & layer_0[1927]; 
    assign out[2387] = layer_0[1845]; 
    assign out[2388] = layer_0[1674] & ~layer_0[1149]; 
    assign out[2389] = ~(layer_0[1991] | layer_0[1767]); 
    assign out[2390] = ~(layer_0[726] | layer_0[83]); 
    assign out[2391] = layer_0[1131] & layer_0[2220]; 
    assign out[2392] = layer_0[1154] | layer_0[1274]; 
    assign out[2393] = ~(layer_0[1073] ^ layer_0[1670]); 
    assign out[2394] = layer_0[1670]; 
    assign out[2395] = ~layer_0[217]; 
    assign out[2396] = ~(layer_0[2047] ^ layer_0[853]); 
    assign out[2397] = layer_0[1611] | layer_0[289]; 
    assign out[2398] = ~(layer_0[2473] ^ layer_0[1054]); 
    assign out[2399] = layer_0[630] ^ layer_0[2276]; 
    assign out[2400] = ~(layer_0[891] ^ layer_0[1420]); 
    assign out[2401] = layer_0[829] ^ layer_0[1852]; 
    assign out[2402] = layer_0[2475]; 
    assign out[2403] = layer_0[2314]; 
    assign out[2404] = ~(layer_0[174] ^ layer_0[1430]); 
    assign out[2405] = ~(layer_0[2526] ^ layer_0[2095]); 
    assign out[2406] = ~layer_0[1473]; 
    assign out[2407] = ~layer_0[1983]; 
    assign out[2408] = layer_0[326] ^ layer_0[717]; 
    assign out[2409] = ~layer_0[469]; 
    assign out[2410] = layer_0[2278] ^ layer_0[610]; 
    assign out[2411] = ~(layer_0[1395] & layer_0[1303]); 
    assign out[2412] = layer_0[670] & ~layer_0[2078]; 
    assign out[2413] = layer_0[2379] ^ layer_0[2121]; 
    assign out[2414] = ~(layer_0[2542] & layer_0[1690]); 
    assign out[2415] = ~layer_0[805]; 
    assign out[2416] = ~(layer_0[967] & layer_0[423]); 
    assign out[2417] = layer_0[1777]; 
    assign out[2418] = layer_0[1293] ^ layer_0[2291]; 
    assign out[2419] = layer_0[2185]; 
    assign out[2420] = layer_0[2404] & ~layer_0[198]; 
    assign out[2421] = ~(layer_0[955] | layer_0[1809]); 
    assign out[2422] = ~(layer_0[1334] ^ layer_0[1071]); 
    assign out[2423] = ~(layer_0[1830] ^ layer_0[323]); 
    assign out[2424] = layer_0[1732] & ~layer_0[903]; 
    assign out[2425] = layer_0[1092]; 
    assign out[2426] = ~layer_0[1861]; 
    assign out[2427] = ~(layer_0[1408] | layer_0[1285]); 
    assign out[2428] = layer_0[228] & ~layer_0[1290]; 
    assign out[2429] = layer_0[2037]; 
    assign out[2430] = layer_0[429] & ~layer_0[1064]; 
    assign out[2431] = layer_0[2183] & ~layer_0[1190]; 
    assign out[2432] = layer_0[604] & ~layer_0[967]; 
    assign out[2433] = layer_0[2315]; 
    assign out[2434] = layer_0[2362] ^ layer_0[1061]; 
    assign out[2435] = ~(layer_0[944] ^ layer_0[2520]); 
    assign out[2436] = layer_0[2247] & ~layer_0[1482]; 
    assign out[2437] = ~(layer_0[2509] ^ layer_0[2215]); 
    assign out[2438] = ~layer_0[1022]; 
    assign out[2439] = layer_0[2075] ^ layer_0[589]; 
    assign out[2440] = ~(layer_0[511] & layer_0[315]); 
    assign out[2441] = ~layer_0[348] | (layer_0[111] & layer_0[348]); 
    assign out[2442] = layer_0[2003]; 
    assign out[2443] = ~layer_0[2542]; 
    assign out[2444] = layer_0[299] ^ layer_0[817]; 
    assign out[2445] = ~(layer_0[1032] ^ layer_0[637]); 
    assign out[2446] = layer_0[227] ^ layer_0[1697]; 
    assign out[2447] = layer_0[311] ^ layer_0[810]; 
    assign out[2448] = ~(layer_0[731] ^ layer_0[1972]); 
    assign out[2449] = ~layer_0[2513] | (layer_0[2513] & layer_0[1506]); 
    assign out[2450] = ~(layer_0[419] ^ layer_0[171]); 
    assign out[2451] = ~layer_0[2224]; 
    assign out[2452] = layer_0[1921]; 
    assign out[2453] = layer_0[1264] ^ layer_0[2310]; 
    assign out[2454] = layer_0[2344] ^ layer_0[1027]; 
    assign out[2455] = layer_0[1534] & ~layer_0[1473]; 
    assign out[2456] = layer_0[388]; 
    assign out[2457] = layer_0[2278] & ~layer_0[1178]; 
    assign out[2458] = layer_0[2083]; 
    assign out[2459] = ~(layer_0[1515] | layer_0[2187]); 
    assign out[2460] = ~layer_0[1805]; 
    assign out[2461] = ~(layer_0[1785] ^ layer_0[1722]); 
    assign out[2462] = layer_0[1575] ^ layer_0[944]; 
    assign out[2463] = ~(layer_0[18] | layer_0[764]); 
    assign out[2464] = layer_0[1206]; 
    assign out[2465] = ~layer_0[1337] | (layer_0[279] & layer_0[1337]); 
    assign out[2466] = ~layer_0[347] | (layer_0[1092] & layer_0[347]); 
    assign out[2467] = ~(layer_0[85] ^ layer_0[261]); 
    assign out[2468] = layer_0[41] & layer_0[2074]; 
    assign out[2469] = layer_0[2545] ^ layer_0[963]; 
    assign out[2470] = layer_0[2276] & layer_0[2014]; 
    assign out[2471] = layer_0[1681] & layer_0[1698]; 
    assign out[2472] = ~(layer_0[1847] | layer_0[2425]); 
    assign out[2473] = ~(layer_0[1722] ^ layer_0[2045]); 
    assign out[2474] = layer_0[1103] & ~layer_0[945]; 
    assign out[2475] = layer_0[2106] ^ layer_0[2223]; 
    assign out[2476] = layer_0[325] ^ layer_0[1049]; 
    assign out[2477] = layer_0[1459] & layer_0[2083]; 
    assign out[2478] = ~(layer_0[2474] ^ layer_0[1573]); 
    assign out[2479] = ~layer_0[2427]; 
    assign out[2480] = ~layer_0[583]; 
    assign out[2481] = layer_0[2503] ^ layer_0[1335]; 
    assign out[2482] = ~layer_0[698]; 
    assign out[2483] = layer_0[1812]; 
    assign out[2484] = ~layer_0[382]; 
    assign out[2485] = layer_0[1964]; 
    assign out[2486] = layer_0[2424]; 
    assign out[2487] = layer_0[2013] & ~layer_0[1786]; 
    assign out[2488] = ~(layer_0[2189] | layer_0[1393]); 
    assign out[2489] = layer_0[1621] & ~layer_0[109]; 
    assign out[2490] = layer_0[2429] & ~layer_0[253]; 
    assign out[2491] = ~layer_0[1923]; 
    assign out[2492] = ~(layer_0[1496] & layer_0[432]); 
    assign out[2493] = ~(layer_0[1925] ^ layer_0[509]); 
    assign out[2494] = layer_0[516] & ~layer_0[197]; 
    assign out[2495] = layer_0[1001] ^ layer_0[449]; 
    assign out[2496] = ~layer_0[682]; 
    assign out[2497] = ~layer_0[1337]; 
    assign out[2498] = ~(layer_0[2517] | layer_0[330]); 
    assign out[2499] = ~(layer_0[2194] ^ layer_0[2509]); 
    assign out[2500] = layer_0[1429] & layer_0[809]; 
    assign out[2501] = ~(layer_0[1010] | layer_0[1727]); 
    assign out[2502] = layer_0[1438] & ~layer_0[2125]; 
    assign out[2503] = ~layer_0[805]; 
    assign out[2504] = ~(layer_0[2201] ^ layer_0[1728]); 
    assign out[2505] = ~layer_0[125]; 
    assign out[2506] = layer_0[1724] ^ layer_0[2235]; 
    assign out[2507] = layer_0[1713] | layer_0[2403]; 
    assign out[2508] = ~layer_0[2425]; 
    assign out[2509] = ~(layer_0[378] ^ layer_0[251]); 
    assign out[2510] = ~layer_0[2336]; 
    assign out[2511] = ~layer_0[201]; 
    assign out[2512] = ~layer_0[2486]; 
    assign out[2513] = ~layer_0[211]; 
    assign out[2514] = layer_0[1721] & layer_0[246]; 
    assign out[2515] = layer_0[1822] & layer_0[2314]; 
    assign out[2516] = ~(layer_0[293] ^ layer_0[155]); 
    assign out[2517] = ~(layer_0[725] | layer_0[2297]); 
    assign out[2518] = layer_0[2335] & ~layer_0[1174]; 
    assign out[2519] = layer_0[815] & ~layer_0[2078]; 
    assign out[2520] = layer_0[1781]; 
    assign out[2521] = layer_0[1162] & layer_0[1030]; 
    assign out[2522] = ~(layer_0[1259] ^ layer_0[805]); 
    assign out[2523] = layer_0[140]; 
    assign out[2524] = ~(layer_0[1955] ^ layer_0[1660]); 
    assign out[2525] = ~(layer_0[1464] ^ layer_0[1359]); 
    assign out[2526] = layer_0[2524] | layer_0[1199]; 
    assign out[2527] = ~layer_0[680]; 
    assign out[2528] = ~(layer_0[611] & layer_0[988]); 
    assign out[2529] = ~layer_0[2079]; 
    assign out[2530] = ~(layer_0[2100] ^ layer_0[101]); 
    assign out[2531] = ~layer_0[1010]; 
    assign out[2532] = ~(layer_0[2350] ^ layer_0[521]); 
    assign out[2533] = ~(layer_0[454] ^ layer_0[637]); 
    assign out[2534] = ~(layer_0[410] ^ layer_0[226]); 
    assign out[2535] = layer_0[2237] | layer_0[2307]; 
    assign out[2536] = ~(layer_0[439] | layer_0[211]); 
    assign out[2537] = layer_0[936] ^ layer_0[233]; 
    assign out[2538] = ~(layer_0[1455] ^ layer_0[1591]); 
    assign out[2539] = ~layer_0[666]; 
    assign out[2540] = layer_0[900]; 
    assign out[2541] = layer_0[971] | layer_0[55]; 
    assign out[2542] = ~(layer_0[33] | layer_0[1334]); 
    assign out[2543] = ~layer_0[913]; 
    assign out[2544] = layer_0[2290] ^ layer_0[1503]; 
    assign out[2545] = ~layer_0[794]; 
    assign out[2546] = layer_0[2532] & ~layer_0[428]; 
    assign out[2547] = layer_0[1085] ^ layer_0[988]; 
    assign out[2548] = ~(layer_0[2032] & layer_0[801]); 
    assign out[2549] = ~(layer_0[1650] & layer_0[198]); 
    assign out[2550] = 1'b0; 
    assign out[2551] = 1'b0; 
    assign out[2552] = 1'b0; 
    assign out[2553] = 1'b0; 
    assign out[2554] = 1'b0; 
    assign out[2555] = 1'b0; 
    assign out[2556] = 1'b0; 
    assign out[2557] = 1'b0; 
    assign out[2558] = 1'b0; 
    assign out[2559] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[254:0] = out[254:0];
    assign categories[509:255] = out[510:256];
    assign categories[764:510] = out[766:512];
    assign categories[1019:765] = out[1022:768];
    assign categories[1274:1020] = out[1278:1024];
    assign categories[1529:1275] = out[1534:1280];
    assign categories[1784:1530] = out[1790:1536];
    assign categories[2039:1785] = out[2046:1792];
    assign categories[2294:2040] = out[2302:2048];
    assign categories[2549:2295] = out[2558:2304];

endmodule
