magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -286 -300 286 300
<< nmos >>
rect -100 -100 100 100
<< ndiff >>
rect -158 85 -100 100
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -100 -100 -85
rect 100 85 158 100
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -100 158 -85
<< ndiffc >>
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
<< psubdiff >>
rect -260 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 260 274
rect -260 153 -226 240
rect -260 85 -226 119
rect 226 153 260 240
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect -260 -240 -226 -153
rect 226 -119 260 -85
rect 226 -240 260 -153
rect -260 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 260 -240
<< psubdiffcont >>
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect -260 119 -226 153
rect 226 119 260 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect -260 -153 -226 -119
rect 226 -153 260 -119
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
<< poly >>
rect -100 172 100 188
rect -100 138 -51 172
rect -17 138 17 172
rect 51 138 100 172
rect -100 100 100 138
rect -100 -138 100 -100
rect -100 -172 -51 -138
rect -17 -172 17 -138
rect 51 -172 100 -138
rect -100 -188 100 -172
<< polycont >>
rect -51 138 -17 172
rect 17 138 51 172
rect -51 -172 -17 -138
rect 17 -172 51 -138
<< locali >>
rect -260 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 260 274
rect -260 153 -226 240
rect -100 138 -53 172
rect -17 138 17 172
rect 53 138 100 172
rect 226 153 260 240
rect -260 85 -226 119
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect -146 85 -112 104
rect -146 17 -112 19
rect -146 -19 -112 -17
rect -146 -104 -112 -85
rect 112 85 146 104
rect 112 17 146 19
rect 112 -19 146 -17
rect 112 -104 146 -85
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect -260 -240 -226 -153
rect -100 -172 -53 -138
rect -17 -172 17 -138
rect 53 -172 100 -138
rect 226 -240 260 -153
rect -260 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 260 -240
<< viali >>
rect -53 138 -51 172
rect -51 138 -19 172
rect 19 138 51 172
rect 51 138 53 172
rect -146 51 -112 53
rect -146 19 -112 51
rect -146 -51 -112 -19
rect -146 -53 -112 -51
rect 112 51 146 53
rect 112 19 146 51
rect 112 -51 146 -19
rect 112 -53 146 -51
rect -53 -172 -51 -138
rect -51 -172 -19 -138
rect 19 -172 51 -138
rect 51 -172 53 -138
<< metal1 >>
rect -96 172 96 178
rect -96 138 -53 172
rect -19 138 19 172
rect 53 138 96 172
rect -96 132 96 138
rect -152 53 -106 100
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -100 -106 -53
rect 106 53 152 100
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -100 152 -53
rect -96 -138 96 -132
rect -96 -172 -53 -138
rect -19 -172 19 -138
rect 53 -172 96 -138
rect -96 -178 96 -172
<< properties >>
string FIXED_BBOX -242 -256 242 256
<< end >>
