magic
tech sky130A
timestamp 1756992108
<< error_p >>
rect -62 140 -33 143
rect 33 140 62 143
rect -62 123 -56 140
rect 33 123 39 140
rect -62 120 -33 123
rect 33 120 62 123
rect -110 -123 -81 -120
rect -14 -123 14 -120
rect 81 -123 110 -120
rect -110 -140 -104 -123
rect -14 -140 -8 -123
rect 81 -140 87 -123
rect -110 -143 -81 -140
rect -14 -143 14 -140
rect 81 -143 110 -140
<< nwell >>
rect -203 -209 203 209
<< pmos >>
rect -103 -100 -88 100
rect -55 -100 -40 100
rect -7 -100 7 100
rect 40 -100 55 100
rect 88 -100 103 100
<< pdiff >>
rect -134 93 -103 100
rect -134 76 -128 93
rect -111 76 -103 93
rect -134 59 -103 76
rect -134 42 -128 59
rect -111 42 -103 59
rect -134 25 -103 42
rect -134 8 -128 25
rect -111 8 -103 25
rect -134 -8 -103 8
rect -134 -25 -128 -8
rect -111 -25 -103 -8
rect -134 -42 -103 -25
rect -134 -59 -128 -42
rect -111 -59 -103 -42
rect -134 -76 -103 -59
rect -134 -93 -128 -76
rect -111 -93 -103 -76
rect -134 -100 -103 -93
rect -88 93 -55 100
rect -88 76 -80 93
rect -63 76 -55 93
rect -88 59 -55 76
rect -88 42 -80 59
rect -63 42 -55 59
rect -88 25 -55 42
rect -88 8 -80 25
rect -63 8 -55 25
rect -88 -8 -55 8
rect -88 -25 -80 -8
rect -63 -25 -55 -8
rect -88 -42 -55 -25
rect -88 -59 -80 -42
rect -63 -59 -55 -42
rect -88 -76 -55 -59
rect -88 -93 -80 -76
rect -63 -93 -55 -76
rect -88 -100 -55 -93
rect -40 93 -7 100
rect -40 76 -32 93
rect -15 76 -7 93
rect -40 59 -7 76
rect -40 42 -32 59
rect -15 42 -7 59
rect -40 25 -7 42
rect -40 8 -32 25
rect -15 8 -7 25
rect -40 -8 -7 8
rect -40 -25 -32 -8
rect -15 -25 -7 -8
rect -40 -42 -7 -25
rect -40 -59 -32 -42
rect -15 -59 -7 -42
rect -40 -76 -7 -59
rect -40 -93 -32 -76
rect -15 -93 -7 -76
rect -40 -100 -7 -93
rect 7 93 40 100
rect 7 76 15 93
rect 32 76 40 93
rect 7 59 40 76
rect 7 42 15 59
rect 32 42 40 59
rect 7 25 40 42
rect 7 8 15 25
rect 32 8 40 25
rect 7 -8 40 8
rect 7 -25 15 -8
rect 32 -25 40 -8
rect 7 -42 40 -25
rect 7 -59 15 -42
rect 32 -59 40 -42
rect 7 -76 40 -59
rect 7 -93 15 -76
rect 32 -93 40 -76
rect 7 -100 40 -93
rect 55 93 88 100
rect 55 76 63 93
rect 80 76 88 93
rect 55 59 88 76
rect 55 42 63 59
rect 80 42 88 59
rect 55 25 88 42
rect 55 8 63 25
rect 80 8 88 25
rect 55 -8 88 8
rect 55 -25 63 -8
rect 80 -25 88 -8
rect 55 -42 88 -25
rect 55 -59 63 -42
rect 80 -59 88 -42
rect 55 -76 88 -59
rect 55 -93 63 -76
rect 80 -93 88 -76
rect 55 -100 88 -93
rect 103 93 134 100
rect 103 76 111 93
rect 128 76 134 93
rect 103 59 134 76
rect 103 42 111 59
rect 128 42 134 59
rect 103 25 134 42
rect 103 8 111 25
rect 128 8 134 25
rect 103 -8 134 8
rect 103 -25 111 -8
rect 128 -25 134 -8
rect 103 -42 134 -25
rect 103 -59 111 -42
rect 128 -59 134 -42
rect 103 -76 134 -59
rect 103 -93 111 -76
rect 128 -93 134 -76
rect 103 -100 134 -93
<< pdiffc >>
rect -128 76 -111 93
rect -128 42 -111 59
rect -128 8 -111 25
rect -128 -25 -111 -8
rect -128 -59 -111 -42
rect -128 -93 -111 -76
rect -80 76 -63 93
rect -80 42 -63 59
rect -80 8 -63 25
rect -80 -25 -63 -8
rect -80 -59 -63 -42
rect -80 -93 -63 -76
rect -32 76 -15 93
rect -32 42 -15 59
rect -32 8 -15 25
rect -32 -25 -15 -8
rect -32 -59 -15 -42
rect -32 -93 -15 -76
rect 15 76 32 93
rect 15 42 32 59
rect 15 8 32 25
rect 15 -25 32 -8
rect 15 -59 32 -42
rect 15 -93 32 -76
rect 63 76 80 93
rect 63 42 80 59
rect 63 8 80 25
rect 63 -25 80 -8
rect 63 -59 80 -42
rect 63 -93 80 -76
rect 111 76 128 93
rect 111 42 128 59
rect 111 8 128 25
rect 111 -25 128 -8
rect 111 -59 128 -42
rect 111 -93 128 -76
<< nsubdiff >>
rect -185 174 -127 191
rect -110 174 -93 191
rect -76 174 -59 191
rect -42 174 -25 191
rect -8 174 8 191
rect 25 174 42 191
rect 59 174 76 191
rect 93 174 110 191
rect 127 174 185 191
rect -185 127 -168 174
rect 168 127 185 174
rect -185 93 -168 110
rect -185 59 -168 76
rect -185 25 -168 42
rect -185 -8 -168 8
rect -185 -42 -168 -25
rect -185 -76 -168 -59
rect -185 -110 -168 -93
rect 168 93 185 110
rect 168 59 185 76
rect 168 25 185 42
rect 168 -8 185 8
rect 168 -42 185 -25
rect 168 -76 185 -59
rect 168 -110 185 -93
rect -185 -174 -168 -127
rect 168 -174 185 -127
rect -185 -191 -127 -174
rect -110 -191 -93 -174
rect -76 -191 -59 -174
rect -42 -191 -25 -174
rect -8 -191 8 -174
rect 25 -191 42 -174
rect 59 -191 76 -174
rect 93 -191 110 -174
rect 127 -191 185 -174
<< nsubdiffcont >>
rect -127 174 -110 191
rect -93 174 -76 191
rect -59 174 -42 191
rect -25 174 -8 191
rect 8 174 25 191
rect 42 174 59 191
rect 76 174 93 191
rect 110 174 127 191
rect -185 110 -168 127
rect 168 110 185 127
rect -185 76 -168 93
rect -185 42 -168 59
rect -185 8 -168 25
rect -185 -25 -168 -8
rect -185 -59 -168 -42
rect -185 -93 -168 -76
rect 168 76 185 93
rect 168 42 185 59
rect 168 8 185 25
rect 168 -25 185 -8
rect 168 -59 185 -42
rect 168 -93 185 -76
rect -185 -127 -168 -110
rect 168 -127 185 -110
rect -127 -191 -110 -174
rect -93 -191 -76 -174
rect -59 -191 -42 -174
rect -25 -191 -8 -174
rect 8 -191 25 -174
rect 42 -191 59 -174
rect 76 -191 93 -174
rect 110 -191 127 -174
<< poly >>
rect -64 140 -31 148
rect -64 123 -56 140
rect -39 123 -31 140
rect -64 115 -31 123
rect 31 140 64 148
rect 31 123 39 140
rect 56 123 64 140
rect 31 115 64 123
rect -103 100 -88 113
rect -55 100 -40 115
rect -7 100 7 113
rect 40 100 55 115
rect 88 100 103 113
rect -103 -115 -88 -100
rect -55 -113 -40 -100
rect -7 -115 7 -100
rect 40 -113 55 -100
rect 88 -115 103 -100
rect -112 -123 -79 -115
rect -112 -140 -104 -123
rect -87 -140 -79 -123
rect -112 -148 -79 -140
rect -16 -123 16 -115
rect -16 -140 -8 -123
rect 8 -140 16 -123
rect -16 -148 16 -140
rect 79 -123 112 -115
rect 79 -140 87 -123
rect 104 -140 112 -123
rect 79 -148 112 -140
<< polycont >>
rect -56 123 -39 140
rect 39 123 56 140
rect -104 -140 -87 -123
rect -8 -140 8 -123
rect 87 -140 104 -123
<< locali >>
rect -185 174 -127 191
rect -110 174 -93 191
rect -76 174 -59 191
rect -42 174 -25 191
rect -8 174 8 191
rect 25 174 42 191
rect 59 174 76 191
rect 93 174 110 191
rect 127 174 185 191
rect -185 127 -168 174
rect -64 123 -56 140
rect -39 123 -31 140
rect 31 123 39 140
rect 56 123 64 140
rect 168 127 185 174
rect -185 93 -168 110
rect -185 59 -168 76
rect -185 25 -168 42
rect -185 -8 -168 8
rect -185 -42 -168 -25
rect -185 -76 -168 -59
rect -185 -110 -168 -93
rect -128 93 -111 102
rect -128 59 -111 63
rect -128 25 -111 27
rect -128 -27 -111 -25
rect -128 -63 -111 -59
rect -128 -102 -111 -93
rect -80 93 -63 102
rect -80 59 -63 63
rect -80 25 -63 27
rect -80 -27 -63 -25
rect -80 -63 -63 -59
rect -80 -102 -63 -93
rect -32 93 -15 102
rect -32 59 -15 63
rect -32 25 -15 27
rect -32 -27 -15 -25
rect -32 -63 -15 -59
rect -32 -102 -15 -93
rect 15 93 32 102
rect 15 59 32 63
rect 15 25 32 27
rect 15 -27 32 -25
rect 15 -63 32 -59
rect 15 -102 32 -93
rect 63 93 80 102
rect 63 59 80 63
rect 63 25 80 27
rect 63 -27 80 -25
rect 63 -63 80 -59
rect 63 -102 80 -93
rect 111 93 128 102
rect 111 59 128 63
rect 111 25 128 27
rect 111 -27 128 -25
rect 111 -63 128 -59
rect 111 -102 128 -93
rect 168 93 185 110
rect 168 59 185 76
rect 168 25 185 42
rect 168 -8 185 8
rect 168 -42 185 -25
rect 168 -76 185 -59
rect 168 -110 185 -93
rect -185 -174 -168 -127
rect -112 -140 -104 -123
rect -87 -140 -79 -123
rect -16 -140 -8 -123
rect 8 -140 16 -123
rect 79 -140 87 -123
rect 104 -140 112 -123
rect 168 -174 185 -127
rect -185 -191 -127 -174
rect -110 -191 -93 -174
rect -76 -191 -59 -174
rect -42 -191 -25 -174
rect -8 -191 8 -174
rect 25 -191 42 -174
rect 59 -191 76 -174
rect 93 -191 110 -174
rect 127 -191 185 -174
<< viali >>
rect -56 123 -39 140
rect 39 123 56 140
rect -128 76 -111 80
rect -128 63 -111 76
rect -128 42 -111 44
rect -128 27 -111 42
rect -128 -8 -111 8
rect -128 -42 -111 -27
rect -128 -44 -111 -42
rect -128 -76 -111 -63
rect -128 -80 -111 -76
rect -80 76 -63 80
rect -80 63 -63 76
rect -80 42 -63 44
rect -80 27 -63 42
rect -80 -8 -63 8
rect -80 -42 -63 -27
rect -80 -44 -63 -42
rect -80 -76 -63 -63
rect -80 -80 -63 -76
rect -32 76 -15 80
rect -32 63 -15 76
rect -32 42 -15 44
rect -32 27 -15 42
rect -32 -8 -15 8
rect -32 -42 -15 -27
rect -32 -44 -15 -42
rect -32 -76 -15 -63
rect -32 -80 -15 -76
rect 15 76 32 80
rect 15 63 32 76
rect 15 42 32 44
rect 15 27 32 42
rect 15 -8 32 8
rect 15 -42 32 -27
rect 15 -44 32 -42
rect 15 -76 32 -63
rect 15 -80 32 -76
rect 63 76 80 80
rect 63 63 80 76
rect 63 42 80 44
rect 63 27 80 42
rect 63 -8 80 8
rect 63 -42 80 -27
rect 63 -44 80 -42
rect 63 -76 80 -63
rect 63 -80 80 -76
rect 111 76 128 80
rect 111 63 128 76
rect 111 42 128 44
rect 111 27 128 42
rect 111 -8 128 8
rect 111 -42 128 -27
rect 111 -44 128 -42
rect 111 -76 128 -63
rect 111 -80 128 -76
rect -104 -140 -87 -123
rect -8 -140 8 -123
rect 87 -140 104 -123
<< metal1 >>
rect -62 140 -33 143
rect -62 123 -56 140
rect -39 123 -33 140
rect -62 120 -33 123
rect 33 140 62 143
rect 33 123 39 140
rect 56 123 62 140
rect 33 120 62 123
rect -131 80 -108 100
rect -131 63 -128 80
rect -111 63 -108 80
rect -131 44 -108 63
rect -131 27 -128 44
rect -111 27 -108 44
rect -131 8 -108 27
rect -131 -8 -128 8
rect -111 -8 -108 8
rect -131 -27 -108 -8
rect -131 -44 -128 -27
rect -111 -44 -108 -27
rect -131 -63 -108 -44
rect -131 -80 -128 -63
rect -111 -80 -108 -63
rect -131 -100 -108 -80
rect -83 80 -60 100
rect -83 63 -80 80
rect -63 63 -60 80
rect -83 44 -60 63
rect -83 27 -80 44
rect -63 27 -60 44
rect -83 8 -60 27
rect -83 -8 -80 8
rect -63 -8 -60 8
rect -83 -27 -60 -8
rect -83 -44 -80 -27
rect -63 -44 -60 -27
rect -83 -63 -60 -44
rect -83 -80 -80 -63
rect -63 -80 -60 -63
rect -83 -100 -60 -80
rect -35 80 -12 100
rect -35 63 -32 80
rect -15 63 -12 80
rect -35 44 -12 63
rect -35 27 -32 44
rect -15 27 -12 44
rect -35 8 -12 27
rect -35 -8 -32 8
rect -15 -8 -12 8
rect -35 -27 -12 -8
rect -35 -44 -32 -27
rect -15 -44 -12 -27
rect -35 -63 -12 -44
rect -35 -80 -32 -63
rect -15 -80 -12 -63
rect -35 -100 -12 -80
rect 12 80 35 100
rect 12 63 15 80
rect 32 63 35 80
rect 12 44 35 63
rect 12 27 15 44
rect 32 27 35 44
rect 12 8 35 27
rect 12 -8 15 8
rect 32 -8 35 8
rect 12 -27 35 -8
rect 12 -44 15 -27
rect 32 -44 35 -27
rect 12 -63 35 -44
rect 12 -80 15 -63
rect 32 -80 35 -63
rect 12 -100 35 -80
rect 60 80 83 100
rect 60 63 63 80
rect 80 63 83 80
rect 60 44 83 63
rect 60 27 63 44
rect 80 27 83 44
rect 60 8 83 27
rect 60 -8 63 8
rect 80 -8 83 8
rect 60 -27 83 -8
rect 60 -44 63 -27
rect 80 -44 83 -27
rect 60 -63 83 -44
rect 60 -80 63 -63
rect 80 -80 83 -63
rect 60 -100 83 -80
rect 108 80 131 100
rect 108 63 111 80
rect 128 63 131 80
rect 108 44 131 63
rect 108 27 111 44
rect 128 27 131 44
rect 108 8 131 27
rect 108 -8 111 8
rect 128 -8 131 8
rect 108 -27 131 -8
rect 108 -44 111 -27
rect 128 -44 131 -27
rect 108 -63 131 -44
rect 108 -80 111 -63
rect 128 -80 131 -63
rect 108 -100 131 -80
rect -110 -123 -81 -120
rect -110 -140 -104 -123
rect -87 -140 -81 -123
rect -110 -143 -81 -140
rect -14 -123 14 -120
rect -14 -140 -8 -123
rect 8 -140 14 -123
rect -14 -143 14 -140
rect 81 -123 110 -120
rect 81 -140 87 -123
rect 104 -140 110 -123
rect 81 -143 110 -140
<< properties >>
string FIXED_BBOX -177 -183 177 183
<< end >>
