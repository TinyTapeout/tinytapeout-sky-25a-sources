magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 512 240
<< ntap >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 464 20 560 60
rect -48 60 560 100
rect -48 100 560 140
rect -48 140 560 180
<< locali >>
rect -48 -20 48 20
rect 464 -20 560 20
rect -48 20 48 60
rect 464 20 560 60
rect -48 60 560 100
rect -48 100 560 140
rect -48 140 560 180
<< ntapc >>
rect 80 100 432 140
<< nwell >>
rect -92 -64 604 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 512 240
<< end >>
