magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -562 -684 562 684
<< pmos >>
rect -366 -464 -266 536
rect -208 -464 -108 536
rect -50 -464 50 536
rect 108 -464 208 536
rect 266 -464 366 536
<< pdiff >>
rect -424 495 -366 536
rect -424 461 -412 495
rect -378 461 -366 495
rect -424 427 -366 461
rect -424 393 -412 427
rect -378 393 -366 427
rect -424 359 -366 393
rect -424 325 -412 359
rect -378 325 -366 359
rect -424 291 -366 325
rect -424 257 -412 291
rect -378 257 -366 291
rect -424 223 -366 257
rect -424 189 -412 223
rect -378 189 -366 223
rect -424 155 -366 189
rect -424 121 -412 155
rect -378 121 -366 155
rect -424 87 -366 121
rect -424 53 -412 87
rect -378 53 -366 87
rect -424 19 -366 53
rect -424 -15 -412 19
rect -378 -15 -366 19
rect -424 -49 -366 -15
rect -424 -83 -412 -49
rect -378 -83 -366 -49
rect -424 -117 -366 -83
rect -424 -151 -412 -117
rect -378 -151 -366 -117
rect -424 -185 -366 -151
rect -424 -219 -412 -185
rect -378 -219 -366 -185
rect -424 -253 -366 -219
rect -424 -287 -412 -253
rect -378 -287 -366 -253
rect -424 -321 -366 -287
rect -424 -355 -412 -321
rect -378 -355 -366 -321
rect -424 -389 -366 -355
rect -424 -423 -412 -389
rect -378 -423 -366 -389
rect -424 -464 -366 -423
rect -266 495 -208 536
rect -266 461 -254 495
rect -220 461 -208 495
rect -266 427 -208 461
rect -266 393 -254 427
rect -220 393 -208 427
rect -266 359 -208 393
rect -266 325 -254 359
rect -220 325 -208 359
rect -266 291 -208 325
rect -266 257 -254 291
rect -220 257 -208 291
rect -266 223 -208 257
rect -266 189 -254 223
rect -220 189 -208 223
rect -266 155 -208 189
rect -266 121 -254 155
rect -220 121 -208 155
rect -266 87 -208 121
rect -266 53 -254 87
rect -220 53 -208 87
rect -266 19 -208 53
rect -266 -15 -254 19
rect -220 -15 -208 19
rect -266 -49 -208 -15
rect -266 -83 -254 -49
rect -220 -83 -208 -49
rect -266 -117 -208 -83
rect -266 -151 -254 -117
rect -220 -151 -208 -117
rect -266 -185 -208 -151
rect -266 -219 -254 -185
rect -220 -219 -208 -185
rect -266 -253 -208 -219
rect -266 -287 -254 -253
rect -220 -287 -208 -253
rect -266 -321 -208 -287
rect -266 -355 -254 -321
rect -220 -355 -208 -321
rect -266 -389 -208 -355
rect -266 -423 -254 -389
rect -220 -423 -208 -389
rect -266 -464 -208 -423
rect -108 495 -50 536
rect -108 461 -96 495
rect -62 461 -50 495
rect -108 427 -50 461
rect -108 393 -96 427
rect -62 393 -50 427
rect -108 359 -50 393
rect -108 325 -96 359
rect -62 325 -50 359
rect -108 291 -50 325
rect -108 257 -96 291
rect -62 257 -50 291
rect -108 223 -50 257
rect -108 189 -96 223
rect -62 189 -50 223
rect -108 155 -50 189
rect -108 121 -96 155
rect -62 121 -50 155
rect -108 87 -50 121
rect -108 53 -96 87
rect -62 53 -50 87
rect -108 19 -50 53
rect -108 -15 -96 19
rect -62 -15 -50 19
rect -108 -49 -50 -15
rect -108 -83 -96 -49
rect -62 -83 -50 -49
rect -108 -117 -50 -83
rect -108 -151 -96 -117
rect -62 -151 -50 -117
rect -108 -185 -50 -151
rect -108 -219 -96 -185
rect -62 -219 -50 -185
rect -108 -253 -50 -219
rect -108 -287 -96 -253
rect -62 -287 -50 -253
rect -108 -321 -50 -287
rect -108 -355 -96 -321
rect -62 -355 -50 -321
rect -108 -389 -50 -355
rect -108 -423 -96 -389
rect -62 -423 -50 -389
rect -108 -464 -50 -423
rect 50 495 108 536
rect 50 461 62 495
rect 96 461 108 495
rect 50 427 108 461
rect 50 393 62 427
rect 96 393 108 427
rect 50 359 108 393
rect 50 325 62 359
rect 96 325 108 359
rect 50 291 108 325
rect 50 257 62 291
rect 96 257 108 291
rect 50 223 108 257
rect 50 189 62 223
rect 96 189 108 223
rect 50 155 108 189
rect 50 121 62 155
rect 96 121 108 155
rect 50 87 108 121
rect 50 53 62 87
rect 96 53 108 87
rect 50 19 108 53
rect 50 -15 62 19
rect 96 -15 108 19
rect 50 -49 108 -15
rect 50 -83 62 -49
rect 96 -83 108 -49
rect 50 -117 108 -83
rect 50 -151 62 -117
rect 96 -151 108 -117
rect 50 -185 108 -151
rect 50 -219 62 -185
rect 96 -219 108 -185
rect 50 -253 108 -219
rect 50 -287 62 -253
rect 96 -287 108 -253
rect 50 -321 108 -287
rect 50 -355 62 -321
rect 96 -355 108 -321
rect 50 -389 108 -355
rect 50 -423 62 -389
rect 96 -423 108 -389
rect 50 -464 108 -423
rect 208 495 266 536
rect 208 461 220 495
rect 254 461 266 495
rect 208 427 266 461
rect 208 393 220 427
rect 254 393 266 427
rect 208 359 266 393
rect 208 325 220 359
rect 254 325 266 359
rect 208 291 266 325
rect 208 257 220 291
rect 254 257 266 291
rect 208 223 266 257
rect 208 189 220 223
rect 254 189 266 223
rect 208 155 266 189
rect 208 121 220 155
rect 254 121 266 155
rect 208 87 266 121
rect 208 53 220 87
rect 254 53 266 87
rect 208 19 266 53
rect 208 -15 220 19
rect 254 -15 266 19
rect 208 -49 266 -15
rect 208 -83 220 -49
rect 254 -83 266 -49
rect 208 -117 266 -83
rect 208 -151 220 -117
rect 254 -151 266 -117
rect 208 -185 266 -151
rect 208 -219 220 -185
rect 254 -219 266 -185
rect 208 -253 266 -219
rect 208 -287 220 -253
rect 254 -287 266 -253
rect 208 -321 266 -287
rect 208 -355 220 -321
rect 254 -355 266 -321
rect 208 -389 266 -355
rect 208 -423 220 -389
rect 254 -423 266 -389
rect 208 -464 266 -423
rect 366 495 424 536
rect 366 461 378 495
rect 412 461 424 495
rect 366 427 424 461
rect 366 393 378 427
rect 412 393 424 427
rect 366 359 424 393
rect 366 325 378 359
rect 412 325 424 359
rect 366 291 424 325
rect 366 257 378 291
rect 412 257 424 291
rect 366 223 424 257
rect 366 189 378 223
rect 412 189 424 223
rect 366 155 424 189
rect 366 121 378 155
rect 412 121 424 155
rect 366 87 424 121
rect 366 53 378 87
rect 412 53 424 87
rect 366 19 424 53
rect 366 -15 378 19
rect 412 -15 424 19
rect 366 -49 424 -15
rect 366 -83 378 -49
rect 412 -83 424 -49
rect 366 -117 424 -83
rect 366 -151 378 -117
rect 412 -151 424 -117
rect 366 -185 424 -151
rect 366 -219 378 -185
rect 412 -219 424 -185
rect 366 -253 424 -219
rect 366 -287 378 -253
rect 412 -287 424 -253
rect 366 -321 424 -287
rect 366 -355 378 -321
rect 412 -355 424 -321
rect 366 -389 424 -355
rect 366 -423 378 -389
rect 412 -423 424 -389
rect 366 -464 424 -423
<< pdiffc >>
rect -412 461 -378 495
rect -412 393 -378 427
rect -412 325 -378 359
rect -412 257 -378 291
rect -412 189 -378 223
rect -412 121 -378 155
rect -412 53 -378 87
rect -412 -15 -378 19
rect -412 -83 -378 -49
rect -412 -151 -378 -117
rect -412 -219 -378 -185
rect -412 -287 -378 -253
rect -412 -355 -378 -321
rect -412 -423 -378 -389
rect -254 461 -220 495
rect -254 393 -220 427
rect -254 325 -220 359
rect -254 257 -220 291
rect -254 189 -220 223
rect -254 121 -220 155
rect -254 53 -220 87
rect -254 -15 -220 19
rect -254 -83 -220 -49
rect -254 -151 -220 -117
rect -254 -219 -220 -185
rect -254 -287 -220 -253
rect -254 -355 -220 -321
rect -254 -423 -220 -389
rect -96 461 -62 495
rect -96 393 -62 427
rect -96 325 -62 359
rect -96 257 -62 291
rect -96 189 -62 223
rect -96 121 -62 155
rect -96 53 -62 87
rect -96 -15 -62 19
rect -96 -83 -62 -49
rect -96 -151 -62 -117
rect -96 -219 -62 -185
rect -96 -287 -62 -253
rect -96 -355 -62 -321
rect -96 -423 -62 -389
rect 62 461 96 495
rect 62 393 96 427
rect 62 325 96 359
rect 62 257 96 291
rect 62 189 96 223
rect 62 121 96 155
rect 62 53 96 87
rect 62 -15 96 19
rect 62 -83 96 -49
rect 62 -151 96 -117
rect 62 -219 96 -185
rect 62 -287 96 -253
rect 62 -355 96 -321
rect 62 -423 96 -389
rect 220 461 254 495
rect 220 393 254 427
rect 220 325 254 359
rect 220 257 254 291
rect 220 189 254 223
rect 220 121 254 155
rect 220 53 254 87
rect 220 -15 254 19
rect 220 -83 254 -49
rect 220 -151 254 -117
rect 220 -219 254 -185
rect 220 -287 254 -253
rect 220 -355 254 -321
rect 220 -423 254 -389
rect 378 461 412 495
rect 378 393 412 427
rect 378 325 412 359
rect 378 257 412 291
rect 378 189 412 223
rect 378 121 412 155
rect 378 53 412 87
rect 378 -15 412 19
rect 378 -83 412 -49
rect 378 -151 412 -117
rect 378 -219 412 -185
rect 378 -287 412 -253
rect 378 -355 412 -321
rect 378 -423 412 -389
<< nsubdiff >>
rect -526 614 -425 648
rect -391 614 -357 648
rect -323 614 -289 648
rect -255 614 -221 648
rect -187 614 -153 648
rect -119 614 -85 648
rect -51 614 -17 648
rect 17 614 51 648
rect 85 614 119 648
rect 153 614 187 648
rect 221 614 255 648
rect 289 614 323 648
rect 357 614 391 648
rect 425 614 526 648
rect -526 527 -492 614
rect -526 459 -492 493
rect -526 391 -492 425
rect -526 323 -492 357
rect -526 255 -492 289
rect -526 187 -492 221
rect -526 119 -492 153
rect -526 51 -492 85
rect -526 -17 -492 17
rect -526 -85 -492 -51
rect -526 -153 -492 -119
rect -526 -221 -492 -187
rect -526 -289 -492 -255
rect -526 -357 -492 -323
rect -526 -425 -492 -391
rect -526 -493 -492 -459
rect 492 527 526 614
rect 492 459 526 493
rect 492 391 526 425
rect 492 323 526 357
rect 492 255 526 289
rect 492 187 526 221
rect 492 119 526 153
rect 492 51 526 85
rect 492 -17 526 17
rect 492 -85 526 -51
rect 492 -153 526 -119
rect 492 -221 526 -187
rect 492 -289 526 -255
rect 492 -357 526 -323
rect 492 -425 526 -391
rect -526 -614 -492 -527
rect 492 -493 526 -459
rect 492 -614 526 -527
rect -526 -648 -425 -614
rect -391 -648 -357 -614
rect -323 -648 -289 -614
rect -255 -648 -221 -614
rect -187 -648 -153 -614
rect -119 -648 -85 -614
rect -51 -648 -17 -614
rect 17 -648 51 -614
rect 85 -648 119 -614
rect 153 -648 187 -614
rect 221 -648 255 -614
rect 289 -648 323 -614
rect 357 -648 391 -614
rect 425 -648 526 -614
<< nsubdiffcont >>
rect -425 614 -391 648
rect -357 614 -323 648
rect -289 614 -255 648
rect -221 614 -187 648
rect -153 614 -119 648
rect -85 614 -51 648
rect -17 614 17 648
rect 51 614 85 648
rect 119 614 153 648
rect 187 614 221 648
rect 255 614 289 648
rect 323 614 357 648
rect 391 614 425 648
rect -526 493 -492 527
rect -526 425 -492 459
rect -526 357 -492 391
rect -526 289 -492 323
rect -526 221 -492 255
rect -526 153 -492 187
rect -526 85 -492 119
rect -526 17 -492 51
rect -526 -51 -492 -17
rect -526 -119 -492 -85
rect -526 -187 -492 -153
rect -526 -255 -492 -221
rect -526 -323 -492 -289
rect -526 -391 -492 -357
rect -526 -459 -492 -425
rect 492 493 526 527
rect 492 425 526 459
rect 492 357 526 391
rect 492 289 526 323
rect 492 221 526 255
rect 492 153 526 187
rect 492 85 526 119
rect 492 17 526 51
rect 492 -51 526 -17
rect 492 -119 526 -85
rect 492 -187 526 -153
rect 492 -255 526 -221
rect 492 -323 526 -289
rect 492 -391 526 -357
rect 492 -459 526 -425
rect -526 -527 -492 -493
rect 492 -527 526 -493
rect -425 -648 -391 -614
rect -357 -648 -323 -614
rect -289 -648 -255 -614
rect -221 -648 -187 -614
rect -153 -648 -119 -614
rect -85 -648 -51 -614
rect -17 -648 17 -614
rect 51 -648 85 -614
rect 119 -648 153 -614
rect 187 -648 221 -614
rect 255 -648 289 -614
rect 323 -648 357 -614
rect 391 -648 425 -614
<< poly >>
rect -366 536 -266 562
rect -208 536 -108 562
rect -50 536 50 562
rect 108 536 208 562
rect 266 536 366 562
rect -366 -511 -266 -464
rect -366 -545 -333 -511
rect -299 -545 -266 -511
rect -366 -561 -266 -545
rect -208 -511 -108 -464
rect -208 -545 -175 -511
rect -141 -545 -108 -511
rect -208 -561 -108 -545
rect -50 -511 50 -464
rect -50 -545 -17 -511
rect 17 -545 50 -511
rect -50 -561 50 -545
rect 108 -511 208 -464
rect 108 -545 141 -511
rect 175 -545 208 -511
rect 108 -561 208 -545
rect 266 -511 366 -464
rect 266 -545 299 -511
rect 333 -545 366 -511
rect 266 -561 366 -545
<< polycont >>
rect -333 -545 -299 -511
rect -175 -545 -141 -511
rect -17 -545 17 -511
rect 141 -545 175 -511
rect 299 -545 333 -511
<< locali >>
rect -526 614 -425 648
rect -391 614 -357 648
rect -323 614 -289 648
rect -255 614 -221 648
rect -187 614 -153 648
rect -119 614 -85 648
rect -51 614 -17 648
rect 17 614 51 648
rect 85 614 119 648
rect 153 614 187 648
rect 221 614 255 648
rect 289 614 323 648
rect 357 614 391 648
rect 425 614 526 648
rect -526 527 -492 614
rect -526 459 -492 493
rect -526 391 -492 425
rect -526 323 -492 357
rect -526 255 -492 289
rect -526 187 -492 221
rect -526 119 -492 153
rect -526 51 -492 85
rect -526 -17 -492 17
rect -526 -85 -492 -51
rect -526 -153 -492 -119
rect -526 -221 -492 -187
rect -526 -289 -492 -255
rect -526 -357 -492 -323
rect -526 -425 -492 -391
rect -526 -493 -492 -459
rect -412 521 -378 540
rect -412 449 -378 461
rect -412 377 -378 393
rect -412 305 -378 325
rect -412 233 -378 257
rect -412 161 -378 189
rect -412 89 -378 121
rect -412 19 -378 53
rect -412 -49 -378 -17
rect -412 -117 -378 -89
rect -412 -185 -378 -161
rect -412 -253 -378 -233
rect -412 -321 -378 -305
rect -412 -389 -378 -377
rect -412 -468 -378 -449
rect -254 521 -220 540
rect -254 449 -220 461
rect -254 377 -220 393
rect -254 305 -220 325
rect -254 233 -220 257
rect -254 161 -220 189
rect -254 89 -220 121
rect -254 19 -220 53
rect -254 -49 -220 -17
rect -254 -117 -220 -89
rect -254 -185 -220 -161
rect -254 -253 -220 -233
rect -254 -321 -220 -305
rect -254 -389 -220 -377
rect -254 -468 -220 -449
rect -96 521 -62 540
rect -96 449 -62 461
rect -96 377 -62 393
rect -96 305 -62 325
rect -96 233 -62 257
rect -96 161 -62 189
rect -96 89 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -17
rect -96 -117 -62 -89
rect -96 -185 -62 -161
rect -96 -253 -62 -233
rect -96 -321 -62 -305
rect -96 -389 -62 -377
rect -96 -468 -62 -449
rect 62 521 96 540
rect 62 449 96 461
rect 62 377 96 393
rect 62 305 96 325
rect 62 233 96 257
rect 62 161 96 189
rect 62 89 96 121
rect 62 19 96 53
rect 62 -49 96 -17
rect 62 -117 96 -89
rect 62 -185 96 -161
rect 62 -253 96 -233
rect 62 -321 96 -305
rect 62 -389 96 -377
rect 62 -468 96 -449
rect 220 521 254 540
rect 220 449 254 461
rect 220 377 254 393
rect 220 305 254 325
rect 220 233 254 257
rect 220 161 254 189
rect 220 89 254 121
rect 220 19 254 53
rect 220 -49 254 -17
rect 220 -117 254 -89
rect 220 -185 254 -161
rect 220 -253 254 -233
rect 220 -321 254 -305
rect 220 -389 254 -377
rect 220 -468 254 -449
rect 378 521 412 540
rect 378 449 412 461
rect 378 377 412 393
rect 378 305 412 325
rect 378 233 412 257
rect 378 161 412 189
rect 378 89 412 121
rect 378 19 412 53
rect 378 -49 412 -17
rect 378 -117 412 -89
rect 378 -185 412 -161
rect 378 -253 412 -233
rect 378 -321 412 -305
rect 378 -389 412 -377
rect 378 -468 412 -449
rect 492 527 526 614
rect 492 459 526 493
rect 492 391 526 425
rect 492 323 526 357
rect 492 255 526 289
rect 492 187 526 221
rect 492 119 526 153
rect 492 51 526 85
rect 492 -17 526 17
rect 492 -85 526 -51
rect 492 -153 526 -119
rect 492 -221 526 -187
rect 492 -289 526 -255
rect 492 -357 526 -323
rect 492 -425 526 -391
rect 492 -493 526 -459
rect -526 -614 -492 -527
rect -366 -545 -333 -511
rect -299 -545 -266 -511
rect -208 -545 -175 -511
rect -141 -545 -108 -511
rect -50 -545 -17 -511
rect 17 -545 50 -511
rect 108 -545 141 -511
rect 175 -545 208 -511
rect 266 -545 299 -511
rect 333 -545 366 -511
rect 492 -614 526 -527
rect -526 -648 -425 -614
rect -391 -648 -357 -614
rect -323 -648 -289 -614
rect -255 -648 -221 -614
rect -187 -648 -153 -614
rect -119 -648 -85 -614
rect -51 -648 -17 -614
rect 17 -648 51 -614
rect 85 -648 119 -614
rect 153 -648 187 -614
rect 221 -648 255 -614
rect 289 -648 323 -614
rect 357 -648 391 -614
rect 425 -648 526 -614
<< viali >>
rect -412 495 -378 521
rect -412 487 -378 495
rect -412 427 -378 449
rect -412 415 -378 427
rect -412 359 -378 377
rect -412 343 -378 359
rect -412 291 -378 305
rect -412 271 -378 291
rect -412 223 -378 233
rect -412 199 -378 223
rect -412 155 -378 161
rect -412 127 -378 155
rect -412 87 -378 89
rect -412 55 -378 87
rect -412 -15 -378 17
rect -412 -17 -378 -15
rect -412 -83 -378 -55
rect -412 -89 -378 -83
rect -412 -151 -378 -127
rect -412 -161 -378 -151
rect -412 -219 -378 -199
rect -412 -233 -378 -219
rect -412 -287 -378 -271
rect -412 -305 -378 -287
rect -412 -355 -378 -343
rect -412 -377 -378 -355
rect -412 -423 -378 -415
rect -412 -449 -378 -423
rect -254 495 -220 521
rect -254 487 -220 495
rect -254 427 -220 449
rect -254 415 -220 427
rect -254 359 -220 377
rect -254 343 -220 359
rect -254 291 -220 305
rect -254 271 -220 291
rect -254 223 -220 233
rect -254 199 -220 223
rect -254 155 -220 161
rect -254 127 -220 155
rect -254 87 -220 89
rect -254 55 -220 87
rect -254 -15 -220 17
rect -254 -17 -220 -15
rect -254 -83 -220 -55
rect -254 -89 -220 -83
rect -254 -151 -220 -127
rect -254 -161 -220 -151
rect -254 -219 -220 -199
rect -254 -233 -220 -219
rect -254 -287 -220 -271
rect -254 -305 -220 -287
rect -254 -355 -220 -343
rect -254 -377 -220 -355
rect -254 -423 -220 -415
rect -254 -449 -220 -423
rect -96 495 -62 521
rect -96 487 -62 495
rect -96 427 -62 449
rect -96 415 -62 427
rect -96 359 -62 377
rect -96 343 -62 359
rect -96 291 -62 305
rect -96 271 -62 291
rect -96 223 -62 233
rect -96 199 -62 223
rect -96 155 -62 161
rect -96 127 -62 155
rect -96 87 -62 89
rect -96 55 -62 87
rect -96 -15 -62 17
rect -96 -17 -62 -15
rect -96 -83 -62 -55
rect -96 -89 -62 -83
rect -96 -151 -62 -127
rect -96 -161 -62 -151
rect -96 -219 -62 -199
rect -96 -233 -62 -219
rect -96 -287 -62 -271
rect -96 -305 -62 -287
rect -96 -355 -62 -343
rect -96 -377 -62 -355
rect -96 -423 -62 -415
rect -96 -449 -62 -423
rect 62 495 96 521
rect 62 487 96 495
rect 62 427 96 449
rect 62 415 96 427
rect 62 359 96 377
rect 62 343 96 359
rect 62 291 96 305
rect 62 271 96 291
rect 62 223 96 233
rect 62 199 96 223
rect 62 155 96 161
rect 62 127 96 155
rect 62 87 96 89
rect 62 55 96 87
rect 62 -15 96 17
rect 62 -17 96 -15
rect 62 -83 96 -55
rect 62 -89 96 -83
rect 62 -151 96 -127
rect 62 -161 96 -151
rect 62 -219 96 -199
rect 62 -233 96 -219
rect 62 -287 96 -271
rect 62 -305 96 -287
rect 62 -355 96 -343
rect 62 -377 96 -355
rect 62 -423 96 -415
rect 62 -449 96 -423
rect 220 495 254 521
rect 220 487 254 495
rect 220 427 254 449
rect 220 415 254 427
rect 220 359 254 377
rect 220 343 254 359
rect 220 291 254 305
rect 220 271 254 291
rect 220 223 254 233
rect 220 199 254 223
rect 220 155 254 161
rect 220 127 254 155
rect 220 87 254 89
rect 220 55 254 87
rect 220 -15 254 17
rect 220 -17 254 -15
rect 220 -83 254 -55
rect 220 -89 254 -83
rect 220 -151 254 -127
rect 220 -161 254 -151
rect 220 -219 254 -199
rect 220 -233 254 -219
rect 220 -287 254 -271
rect 220 -305 254 -287
rect 220 -355 254 -343
rect 220 -377 254 -355
rect 220 -423 254 -415
rect 220 -449 254 -423
rect 378 495 412 521
rect 378 487 412 495
rect 378 427 412 449
rect 378 415 412 427
rect 378 359 412 377
rect 378 343 412 359
rect 378 291 412 305
rect 378 271 412 291
rect 378 223 412 233
rect 378 199 412 223
rect 378 155 412 161
rect 378 127 412 155
rect 378 87 412 89
rect 378 55 412 87
rect 378 -15 412 17
rect 378 -17 412 -15
rect 378 -83 412 -55
rect 378 -89 412 -83
rect 378 -151 412 -127
rect 378 -161 412 -151
rect 378 -219 412 -199
rect 378 -233 412 -219
rect 378 -287 412 -271
rect 378 -305 412 -287
rect 378 -355 412 -343
rect 378 -377 412 -355
rect 378 -423 412 -415
rect 378 -449 412 -423
rect -333 -545 -299 -511
rect -175 -545 -141 -511
rect -17 -545 17 -511
rect 141 -545 175 -511
rect 299 -545 333 -511
<< metal1 >>
rect -418 521 -372 536
rect -418 487 -412 521
rect -378 487 -372 521
rect -418 449 -372 487
rect -418 415 -412 449
rect -378 415 -372 449
rect -418 377 -372 415
rect -418 343 -412 377
rect -378 343 -372 377
rect -418 305 -372 343
rect -418 271 -412 305
rect -378 271 -372 305
rect -418 233 -372 271
rect -418 199 -412 233
rect -378 199 -372 233
rect -418 161 -372 199
rect -418 127 -412 161
rect -378 127 -372 161
rect -418 89 -372 127
rect -418 55 -412 89
rect -378 55 -372 89
rect -418 17 -372 55
rect -418 -17 -412 17
rect -378 -17 -372 17
rect -418 -55 -372 -17
rect -418 -89 -412 -55
rect -378 -89 -372 -55
rect -418 -127 -372 -89
rect -418 -161 -412 -127
rect -378 -161 -372 -127
rect -418 -199 -372 -161
rect -418 -233 -412 -199
rect -378 -233 -372 -199
rect -418 -271 -372 -233
rect -418 -305 -412 -271
rect -378 -305 -372 -271
rect -418 -343 -372 -305
rect -418 -377 -412 -343
rect -378 -377 -372 -343
rect -418 -415 -372 -377
rect -418 -449 -412 -415
rect -378 -449 -372 -415
rect -418 -464 -372 -449
rect -260 521 -214 536
rect -260 487 -254 521
rect -220 487 -214 521
rect -260 449 -214 487
rect -260 415 -254 449
rect -220 415 -214 449
rect -260 377 -214 415
rect -260 343 -254 377
rect -220 343 -214 377
rect -260 305 -214 343
rect -260 271 -254 305
rect -220 271 -214 305
rect -260 233 -214 271
rect -260 199 -254 233
rect -220 199 -214 233
rect -260 161 -214 199
rect -260 127 -254 161
rect -220 127 -214 161
rect -260 89 -214 127
rect -260 55 -254 89
rect -220 55 -214 89
rect -260 17 -214 55
rect -260 -17 -254 17
rect -220 -17 -214 17
rect -260 -55 -214 -17
rect -260 -89 -254 -55
rect -220 -89 -214 -55
rect -260 -127 -214 -89
rect -260 -161 -254 -127
rect -220 -161 -214 -127
rect -260 -199 -214 -161
rect -260 -233 -254 -199
rect -220 -233 -214 -199
rect -260 -271 -214 -233
rect -260 -305 -254 -271
rect -220 -305 -214 -271
rect -260 -343 -214 -305
rect -260 -377 -254 -343
rect -220 -377 -214 -343
rect -260 -415 -214 -377
rect -260 -449 -254 -415
rect -220 -449 -214 -415
rect -260 -464 -214 -449
rect -102 521 -56 536
rect -102 487 -96 521
rect -62 487 -56 521
rect -102 449 -56 487
rect -102 415 -96 449
rect -62 415 -56 449
rect -102 377 -56 415
rect -102 343 -96 377
rect -62 343 -56 377
rect -102 305 -56 343
rect -102 271 -96 305
rect -62 271 -56 305
rect -102 233 -56 271
rect -102 199 -96 233
rect -62 199 -56 233
rect -102 161 -56 199
rect -102 127 -96 161
rect -62 127 -56 161
rect -102 89 -56 127
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -127 -56 -89
rect -102 -161 -96 -127
rect -62 -161 -56 -127
rect -102 -199 -56 -161
rect -102 -233 -96 -199
rect -62 -233 -56 -199
rect -102 -271 -56 -233
rect -102 -305 -96 -271
rect -62 -305 -56 -271
rect -102 -343 -56 -305
rect -102 -377 -96 -343
rect -62 -377 -56 -343
rect -102 -415 -56 -377
rect -102 -449 -96 -415
rect -62 -449 -56 -415
rect -102 -464 -56 -449
rect 56 521 102 536
rect 56 487 62 521
rect 96 487 102 521
rect 56 449 102 487
rect 56 415 62 449
rect 96 415 102 449
rect 56 377 102 415
rect 56 343 62 377
rect 96 343 102 377
rect 56 305 102 343
rect 56 271 62 305
rect 96 271 102 305
rect 56 233 102 271
rect 56 199 62 233
rect 96 199 102 233
rect 56 161 102 199
rect 56 127 62 161
rect 96 127 102 161
rect 56 89 102 127
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -127 102 -89
rect 56 -161 62 -127
rect 96 -161 102 -127
rect 56 -199 102 -161
rect 56 -233 62 -199
rect 96 -233 102 -199
rect 56 -271 102 -233
rect 56 -305 62 -271
rect 96 -305 102 -271
rect 56 -343 102 -305
rect 56 -377 62 -343
rect 96 -377 102 -343
rect 56 -415 102 -377
rect 56 -449 62 -415
rect 96 -449 102 -415
rect 56 -464 102 -449
rect 214 521 260 536
rect 214 487 220 521
rect 254 487 260 521
rect 214 449 260 487
rect 214 415 220 449
rect 254 415 260 449
rect 214 377 260 415
rect 214 343 220 377
rect 254 343 260 377
rect 214 305 260 343
rect 214 271 220 305
rect 254 271 260 305
rect 214 233 260 271
rect 214 199 220 233
rect 254 199 260 233
rect 214 161 260 199
rect 214 127 220 161
rect 254 127 260 161
rect 214 89 260 127
rect 214 55 220 89
rect 254 55 260 89
rect 214 17 260 55
rect 214 -17 220 17
rect 254 -17 260 17
rect 214 -55 260 -17
rect 214 -89 220 -55
rect 254 -89 260 -55
rect 214 -127 260 -89
rect 214 -161 220 -127
rect 254 -161 260 -127
rect 214 -199 260 -161
rect 214 -233 220 -199
rect 254 -233 260 -199
rect 214 -271 260 -233
rect 214 -305 220 -271
rect 254 -305 260 -271
rect 214 -343 260 -305
rect 214 -377 220 -343
rect 254 -377 260 -343
rect 214 -415 260 -377
rect 214 -449 220 -415
rect 254 -449 260 -415
rect 214 -464 260 -449
rect 372 521 418 536
rect 372 487 378 521
rect 412 487 418 521
rect 372 449 418 487
rect 372 415 378 449
rect 412 415 418 449
rect 372 377 418 415
rect 372 343 378 377
rect 412 343 418 377
rect 372 305 418 343
rect 372 271 378 305
rect 412 271 418 305
rect 372 233 418 271
rect 372 199 378 233
rect 412 199 418 233
rect 372 161 418 199
rect 372 127 378 161
rect 412 127 418 161
rect 372 89 418 127
rect 372 55 378 89
rect 412 55 418 89
rect 372 17 418 55
rect 372 -17 378 17
rect 412 -17 418 17
rect 372 -55 418 -17
rect 372 -89 378 -55
rect 412 -89 418 -55
rect 372 -127 418 -89
rect 372 -161 378 -127
rect 412 -161 418 -127
rect 372 -199 418 -161
rect 372 -233 378 -199
rect 412 -233 418 -199
rect 372 -271 418 -233
rect 372 -305 378 -271
rect 412 -305 418 -271
rect 372 -343 418 -305
rect 372 -377 378 -343
rect 412 -377 418 -343
rect 372 -415 418 -377
rect 372 -449 378 -415
rect 412 -449 418 -415
rect 372 -464 418 -449
rect -362 -511 -270 -505
rect -362 -545 -333 -511
rect -299 -545 -270 -511
rect -362 -551 -270 -545
rect -204 -511 -112 -505
rect -204 -545 -175 -511
rect -141 -545 -112 -511
rect -204 -551 -112 -545
rect -46 -511 46 -505
rect -46 -545 -17 -511
rect 17 -545 46 -511
rect -46 -551 46 -545
rect 112 -511 204 -505
rect 112 -545 141 -511
rect 175 -545 204 -511
rect 112 -551 204 -545
rect 270 -511 362 -505
rect 270 -545 299 -511
rect 333 -545 362 -511
rect 270 -551 362 -545
<< properties >>
string FIXED_BBOX -509 -631 509 631
<< end >>
