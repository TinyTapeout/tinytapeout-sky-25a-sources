magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 1152 1280
use JNWATR_NCH_4CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 576 240
use JNWATR_NCH_4C1F2 xa2 
transform 1 0 0 0 1 240
box 0 240 576 640
use JNWATR_NCH_4C5F0 xa3 
transform 1 0 0 0 1 640
box 0 640 576 1040
use JNWATR_NCH_4CTAPTOP xa4 
transform 1 0 0 0 1 1040
box 0 1040 576 1280
use JNWATR_NCH_4CTAPBOT xb1 
transform 1 0 576 0 1 0
box 576 0 1152 240
use JNWATR_NCH_4C1F2 xb2 
transform 1 0 576 0 1 240
box 576 240 1152 640
use JNWATR_NCH_4C5F0 xb3 
transform 1 0 576 0 1 640
box 576 640 1152 1040
use JNWATR_NCH_4CTAPTOP xb4 
transform 1 0 576 0 1 1040
box 576 1040 1152 1280
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1152 1280
<< end >>
