
*-------------------------------------------------------------
* JNWATR_PCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_2C1F2 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.22  nf=2  w=0.96  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_2CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_2CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_2CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_2CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_2C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_2C5F0 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.94  nf=2  w=0.96  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_2CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_2CTOP 
xa1  JNWATR_PCH_2CTAPBOT
xa2 D2 G2 S2 B JNWATR_PCH_2C1F2
xa3 D3 G3 S3 B JNWATR_PCH_2C5F0
xa4  JNWATR_PCH_2CTAPTOP
xb1  JNWATR_PCH_2CTAPBOT
xb2 D4 G4 S4 B JNWATR_PCH_2C1F2
xb3 D5 G5 S5 B JNWATR_PCH_2C5F0
xb4  JNWATR_PCH_2CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_4C1F2 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.22  nf=2  w=1.6  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_4CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_4CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_4CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_4CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_4C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_4C5F0 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.94  nf=2  w=1.6  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_4CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_4CTOP 
xa1  JNWATR_PCH_4CTAPBOT
xa2 D2 G2 S2 B JNWATR_PCH_4C1F2
xa3 D3 G3 S3 B JNWATR_PCH_4C5F0
xa4  JNWATR_PCH_4CTAPTOP
xb1  JNWATR_PCH_4CTAPBOT
xb2 D4 G4 S4 B JNWATR_PCH_4C1F2
xb3 D5 G5 S5 B JNWATR_PCH_4C5F0
xb4  JNWATR_PCH_4CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_8C1F2 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.22  nf=2  w=2.88  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_8CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_8CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_8CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_8CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_8C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_8C5F0 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.94  nf=2  w=2.88  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_8CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_8CTOP 
xa1  JNWATR_PCH_8CTAPBOT
xa2 D2 G2 S2 B JNWATR_PCH_8C1F2
xa3 D3 G3 S3 B JNWATR_PCH_8C5F0
xa4  JNWATR_PCH_8CTAPTOP
xb1  JNWATR_PCH_8CTAPBOT
xb2 D4 G4 S4 B JNWATR_PCH_8C1F2
xb3 D5 G5 S5 B JNWATR_PCH_8C5F0
xb4  JNWATR_PCH_8CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_12C1F2 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.22  nf=2  w=4.16  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_12CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_12CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_12CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_12CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_12C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_12C5F0 D G S B
M1 D G S B sky130_fd_pr__pfet_01v8  l=0.94  nf=2  w=4.16  
.ENDS

*-------------------------------------------------------------
* JNWATR_PCH_12CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_PCH_12CTOP 
xa1  JNWATR_PCH_12CTAPBOT
xa2 D2 G2 S2 B JNWATR_PCH_12C1F2
xa3 D3 G3 S3 B JNWATR_PCH_12C5F0
xa4  JNWATR_PCH_12CTAPTOP
xb1  JNWATR_PCH_12CTAPBOT
xb2 D4 G4 S4 B JNWATR_PCH_12C1F2
xb3 D5 G5 S5 B JNWATR_PCH_12C5F0
xb4  JNWATR_PCH_12CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_2C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_2C1F2 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.22  nf=2  w=0.96  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_2CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_2CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_2CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_2CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_2C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_2C5F0 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.94  nf=2  w=0.96  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_2CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_2CTOP 
xa1  JNWATR_NCH_2CTAPBOT
xa2 D2 G2 S2 B JNWATR_NCH_2C1F2
xa3 D3 G3 S3 B JNWATR_NCH_2C5F0
xa4  JNWATR_NCH_2CTAPTOP
xb1  JNWATR_NCH_2CTAPBOT
xb2 D4 G4 S4 B JNWATR_NCH_2C1F2
xb3 D5 G5 S5 B JNWATR_NCH_2C5F0
xb4  JNWATR_NCH_2CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_4C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_4C1F2 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.22  nf=2  w=1.6  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_4CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_4CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_4CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_4CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_4C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_4C5F0 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.94  nf=2  w=1.6  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_4CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_4CTOP 
xa1  JNWATR_NCH_4CTAPBOT
xa2 D2 G2 S2 B JNWATR_NCH_4C1F2
xa3 D3 G3 S3 B JNWATR_NCH_4C5F0
xa4  JNWATR_NCH_4CTAPTOP
xb1  JNWATR_NCH_4CTAPBOT
xb2 D4 G4 S4 B JNWATR_NCH_4C1F2
xb3 D5 G5 S5 B JNWATR_NCH_4C5F0
xb4  JNWATR_NCH_4CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_8C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_8C1F2 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.22  nf=2  w=2.88  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_8CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_8CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_8CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_8CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_8C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_8C5F0 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.94  nf=2  w=2.88  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_8CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_8CTOP 
xa1  JNWATR_NCH_8CTAPBOT
xa2 D2 G2 S2 B JNWATR_NCH_8C1F2
xa3 D3 G3 S3 B JNWATR_NCH_8C5F0
xa4  JNWATR_NCH_8CTAPTOP
xb1  JNWATR_NCH_8CTAPBOT
xb2 D4 G4 S4 B JNWATR_NCH_8C1F2
xb3 D5 G5 S5 B JNWATR_NCH_8C5F0
xb4  JNWATR_NCH_8CTAPTOP
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_12C1F2 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_12C1F2 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.22  nf=2  w=4.16  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_12CTAPTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_12CTAPTOP 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_12CTAPBOT <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_12CTAPBOT 
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_12C5F0 <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_12C5F0 D G S B
M1 D G S B sky130_fd_pr__nfet_01v8  l=0.94  nf=2  w=4.16  
.ENDS

*-------------------------------------------------------------
* JNWATR_NCH_12CTOP <class 'cicpy.core.layoutcell.LayoutCell'>
*-------------------------------------------------------------
.SUBCKT JNWATR_NCH_12CTOP 
xa1  JNWATR_NCH_12CTAPBOT
xa2 D2 G2 S2 B JNWATR_NCH_12C1F2
xa3 D3 G3 S3 B JNWATR_NCH_12C5F0
xa4  JNWATR_NCH_12CTAPTOP
xb1  JNWATR_NCH_12CTAPBOT
xb2 D4 G4 S4 B JNWATR_NCH_12C1F2
xb3 D5 G5 S5 B JNWATR_NCH_12C5F0
xb4  JNWATR_NCH_12CTAPTOP
.ENDS
