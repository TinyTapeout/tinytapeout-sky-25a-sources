magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -236 -500 236 500
<< nmos >>
rect -50 -300 50 300
<< ndiff >>
rect -108 255 -50 300
rect -108 221 -96 255
rect -62 221 -50 255
rect -108 187 -50 221
rect -108 153 -96 187
rect -62 153 -50 187
rect -108 119 -50 153
rect -108 85 -96 119
rect -62 85 -50 119
rect -108 51 -50 85
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -85 -50 -51
rect -108 -119 -96 -85
rect -62 -119 -50 -85
rect -108 -153 -50 -119
rect -108 -187 -96 -153
rect -62 -187 -50 -153
rect -108 -221 -50 -187
rect -108 -255 -96 -221
rect -62 -255 -50 -221
rect -108 -300 -50 -255
rect 50 255 108 300
rect 50 221 62 255
rect 96 221 108 255
rect 50 187 108 221
rect 50 153 62 187
rect 96 153 108 187
rect 50 119 108 153
rect 50 85 62 119
rect 96 85 108 119
rect 50 51 108 85
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -85 108 -51
rect 50 -119 62 -85
rect 96 -119 108 -85
rect 50 -153 108 -119
rect 50 -187 62 -153
rect 96 -187 108 -153
rect 50 -221 108 -187
rect 50 -255 62 -221
rect 96 -255 108 -221
rect 50 -300 108 -255
<< ndiffc >>
rect -96 221 -62 255
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect -96 -255 -62 -221
rect 62 221 96 255
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
rect 62 -255 96 -221
<< psubdiff >>
rect -210 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 210 474
rect -210 357 -176 440
rect -210 289 -176 323
rect 176 357 210 440
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect -210 -440 -176 -357
rect 176 -323 210 -289
rect 176 -440 210 -357
rect -210 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 210 -440
<< psubdiffcont >>
rect -85 440 -51 474
rect -17 440 17 474
rect 51 440 85 474
rect -210 323 -176 357
rect 176 323 210 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect -210 -357 -176 -323
rect 176 -357 210 -323
rect -85 -474 -51 -440
rect -17 -474 17 -440
rect 51 -474 85 -440
<< poly >>
rect -50 372 50 388
rect -50 338 -17 372
rect 17 338 50 372
rect -50 300 50 338
rect -50 -338 50 -300
rect -50 -372 -17 -338
rect 17 -372 50 -338
rect -50 -388 50 -372
<< polycont >>
rect -17 338 17 372
rect -17 -372 17 -338
<< locali >>
rect -210 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 210 474
rect -210 357 -176 440
rect -50 338 -17 372
rect 17 338 50 372
rect 176 357 210 440
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -96 269 -62 304
rect -96 197 -62 221
rect -96 125 -62 153
rect -96 53 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -53
rect -96 -153 -62 -125
rect -96 -221 -62 -197
rect -96 -304 -62 -269
rect 62 269 96 304
rect 62 197 96 221
rect 62 125 96 153
rect 62 53 96 85
rect 62 -17 96 17
rect 62 -85 96 -53
rect 62 -153 96 -125
rect 62 -221 96 -197
rect 62 -304 96 -269
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect -210 -440 -176 -357
rect -50 -372 -17 -338
rect 17 -372 50 -338
rect 176 -440 210 -357
rect -210 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 210 -440
<< viali >>
rect -17 338 17 372
rect -96 255 -62 269
rect -96 235 -62 255
rect -96 187 -62 197
rect -96 163 -62 187
rect -96 119 -62 125
rect -96 91 -62 119
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect -96 -119 -62 -91
rect -96 -125 -62 -119
rect -96 -187 -62 -163
rect -96 -197 -62 -187
rect -96 -255 -62 -235
rect -96 -269 -62 -255
rect 62 255 96 269
rect 62 235 96 255
rect 62 187 96 197
rect 62 163 96 187
rect 62 119 96 125
rect 62 91 96 119
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect 62 -119 96 -91
rect 62 -125 96 -119
rect 62 -187 96 -163
rect 62 -197 96 -187
rect 62 -255 96 -235
rect 62 -269 96 -255
rect -17 -372 17 -338
<< metal1 >>
rect -46 372 46 378
rect -46 338 -17 372
rect 17 338 46 372
rect -46 332 46 338
rect -102 269 -56 300
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -300 -56 -269
rect 56 269 102 300
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -300 102 -269
rect -46 -338 46 -332
rect -46 -372 -17 -338
rect 17 -372 46 -338
rect -46 -378 46 -372
<< properties >>
string FIXED_BBOX -192 -456 192 456
<< end >>
