magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 576 240
<< ptap >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 528 20 624 60
rect -48 60 624 100
rect -48 100 624 140
rect -48 140 624 180
<< locali >>
rect -48 -20 48 20
rect 528 -20 624 20
rect -48 20 48 60
rect 528 20 624 60
rect -48 60 624 100
rect -48 100 624 140
rect -48 140 624 180
<< ptapc >>
rect 80 100 496 140
<< pwell >>
rect -92 -64 668 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 576 240
<< end >>
