magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -206 1581 -148 1587
rect -88 1581 -30 1587
rect 30 1581 88 1587
rect 148 1581 206 1587
rect -206 1547 -194 1581
rect -88 1547 -76 1581
rect 30 1547 42 1581
rect 148 1547 160 1581
rect -206 1541 -148 1547
rect -88 1541 -30 1547
rect 30 1541 88 1547
rect 148 1541 206 1547
rect -206 -1547 -148 -1541
rect -88 -1547 -30 -1541
rect 30 -1547 88 -1541
rect 148 -1547 206 -1541
rect -206 -1581 -194 -1547
rect -88 -1581 -76 -1547
rect 30 -1581 42 -1547
rect 148 -1581 160 -1547
rect -206 -1587 -148 -1581
rect -88 -1587 -30 -1581
rect 30 -1587 88 -1581
rect 148 -1587 206 -1581
<< nwell >>
rect -403 -1719 403 1719
<< pmos >>
rect -207 -1500 -147 1500
rect -89 -1500 -29 1500
rect 29 -1500 89 1500
rect 147 -1500 207 1500
<< pdiff >>
rect -265 1479 -207 1500
rect -265 1445 -253 1479
rect -219 1445 -207 1479
rect -265 1411 -207 1445
rect -265 1377 -253 1411
rect -219 1377 -207 1411
rect -265 1343 -207 1377
rect -265 1309 -253 1343
rect -219 1309 -207 1343
rect -265 1275 -207 1309
rect -265 1241 -253 1275
rect -219 1241 -207 1275
rect -265 1207 -207 1241
rect -265 1173 -253 1207
rect -219 1173 -207 1207
rect -265 1139 -207 1173
rect -265 1105 -253 1139
rect -219 1105 -207 1139
rect -265 1071 -207 1105
rect -265 1037 -253 1071
rect -219 1037 -207 1071
rect -265 1003 -207 1037
rect -265 969 -253 1003
rect -219 969 -207 1003
rect -265 935 -207 969
rect -265 901 -253 935
rect -219 901 -207 935
rect -265 867 -207 901
rect -265 833 -253 867
rect -219 833 -207 867
rect -265 799 -207 833
rect -265 765 -253 799
rect -219 765 -207 799
rect -265 731 -207 765
rect -265 697 -253 731
rect -219 697 -207 731
rect -265 663 -207 697
rect -265 629 -253 663
rect -219 629 -207 663
rect -265 595 -207 629
rect -265 561 -253 595
rect -219 561 -207 595
rect -265 527 -207 561
rect -265 493 -253 527
rect -219 493 -207 527
rect -265 459 -207 493
rect -265 425 -253 459
rect -219 425 -207 459
rect -265 391 -207 425
rect -265 357 -253 391
rect -219 357 -207 391
rect -265 323 -207 357
rect -265 289 -253 323
rect -219 289 -207 323
rect -265 255 -207 289
rect -265 221 -253 255
rect -219 221 -207 255
rect -265 187 -207 221
rect -265 153 -253 187
rect -219 153 -207 187
rect -265 119 -207 153
rect -265 85 -253 119
rect -219 85 -207 119
rect -265 51 -207 85
rect -265 17 -253 51
rect -219 17 -207 51
rect -265 -17 -207 17
rect -265 -51 -253 -17
rect -219 -51 -207 -17
rect -265 -85 -207 -51
rect -265 -119 -253 -85
rect -219 -119 -207 -85
rect -265 -153 -207 -119
rect -265 -187 -253 -153
rect -219 -187 -207 -153
rect -265 -221 -207 -187
rect -265 -255 -253 -221
rect -219 -255 -207 -221
rect -265 -289 -207 -255
rect -265 -323 -253 -289
rect -219 -323 -207 -289
rect -265 -357 -207 -323
rect -265 -391 -253 -357
rect -219 -391 -207 -357
rect -265 -425 -207 -391
rect -265 -459 -253 -425
rect -219 -459 -207 -425
rect -265 -493 -207 -459
rect -265 -527 -253 -493
rect -219 -527 -207 -493
rect -265 -561 -207 -527
rect -265 -595 -253 -561
rect -219 -595 -207 -561
rect -265 -629 -207 -595
rect -265 -663 -253 -629
rect -219 -663 -207 -629
rect -265 -697 -207 -663
rect -265 -731 -253 -697
rect -219 -731 -207 -697
rect -265 -765 -207 -731
rect -265 -799 -253 -765
rect -219 -799 -207 -765
rect -265 -833 -207 -799
rect -265 -867 -253 -833
rect -219 -867 -207 -833
rect -265 -901 -207 -867
rect -265 -935 -253 -901
rect -219 -935 -207 -901
rect -265 -969 -207 -935
rect -265 -1003 -253 -969
rect -219 -1003 -207 -969
rect -265 -1037 -207 -1003
rect -265 -1071 -253 -1037
rect -219 -1071 -207 -1037
rect -265 -1105 -207 -1071
rect -265 -1139 -253 -1105
rect -219 -1139 -207 -1105
rect -265 -1173 -207 -1139
rect -265 -1207 -253 -1173
rect -219 -1207 -207 -1173
rect -265 -1241 -207 -1207
rect -265 -1275 -253 -1241
rect -219 -1275 -207 -1241
rect -265 -1309 -207 -1275
rect -265 -1343 -253 -1309
rect -219 -1343 -207 -1309
rect -265 -1377 -207 -1343
rect -265 -1411 -253 -1377
rect -219 -1411 -207 -1377
rect -265 -1445 -207 -1411
rect -265 -1479 -253 -1445
rect -219 -1479 -207 -1445
rect -265 -1500 -207 -1479
rect -147 1479 -89 1500
rect -147 1445 -135 1479
rect -101 1445 -89 1479
rect -147 1411 -89 1445
rect -147 1377 -135 1411
rect -101 1377 -89 1411
rect -147 1343 -89 1377
rect -147 1309 -135 1343
rect -101 1309 -89 1343
rect -147 1275 -89 1309
rect -147 1241 -135 1275
rect -101 1241 -89 1275
rect -147 1207 -89 1241
rect -147 1173 -135 1207
rect -101 1173 -89 1207
rect -147 1139 -89 1173
rect -147 1105 -135 1139
rect -101 1105 -89 1139
rect -147 1071 -89 1105
rect -147 1037 -135 1071
rect -101 1037 -89 1071
rect -147 1003 -89 1037
rect -147 969 -135 1003
rect -101 969 -89 1003
rect -147 935 -89 969
rect -147 901 -135 935
rect -101 901 -89 935
rect -147 867 -89 901
rect -147 833 -135 867
rect -101 833 -89 867
rect -147 799 -89 833
rect -147 765 -135 799
rect -101 765 -89 799
rect -147 731 -89 765
rect -147 697 -135 731
rect -101 697 -89 731
rect -147 663 -89 697
rect -147 629 -135 663
rect -101 629 -89 663
rect -147 595 -89 629
rect -147 561 -135 595
rect -101 561 -89 595
rect -147 527 -89 561
rect -147 493 -135 527
rect -101 493 -89 527
rect -147 459 -89 493
rect -147 425 -135 459
rect -101 425 -89 459
rect -147 391 -89 425
rect -147 357 -135 391
rect -101 357 -89 391
rect -147 323 -89 357
rect -147 289 -135 323
rect -101 289 -89 323
rect -147 255 -89 289
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -289 -89 -255
rect -147 -323 -135 -289
rect -101 -323 -89 -289
rect -147 -357 -89 -323
rect -147 -391 -135 -357
rect -101 -391 -89 -357
rect -147 -425 -89 -391
rect -147 -459 -135 -425
rect -101 -459 -89 -425
rect -147 -493 -89 -459
rect -147 -527 -135 -493
rect -101 -527 -89 -493
rect -147 -561 -89 -527
rect -147 -595 -135 -561
rect -101 -595 -89 -561
rect -147 -629 -89 -595
rect -147 -663 -135 -629
rect -101 -663 -89 -629
rect -147 -697 -89 -663
rect -147 -731 -135 -697
rect -101 -731 -89 -697
rect -147 -765 -89 -731
rect -147 -799 -135 -765
rect -101 -799 -89 -765
rect -147 -833 -89 -799
rect -147 -867 -135 -833
rect -101 -867 -89 -833
rect -147 -901 -89 -867
rect -147 -935 -135 -901
rect -101 -935 -89 -901
rect -147 -969 -89 -935
rect -147 -1003 -135 -969
rect -101 -1003 -89 -969
rect -147 -1037 -89 -1003
rect -147 -1071 -135 -1037
rect -101 -1071 -89 -1037
rect -147 -1105 -89 -1071
rect -147 -1139 -135 -1105
rect -101 -1139 -89 -1105
rect -147 -1173 -89 -1139
rect -147 -1207 -135 -1173
rect -101 -1207 -89 -1173
rect -147 -1241 -89 -1207
rect -147 -1275 -135 -1241
rect -101 -1275 -89 -1241
rect -147 -1309 -89 -1275
rect -147 -1343 -135 -1309
rect -101 -1343 -89 -1309
rect -147 -1377 -89 -1343
rect -147 -1411 -135 -1377
rect -101 -1411 -89 -1377
rect -147 -1445 -89 -1411
rect -147 -1479 -135 -1445
rect -101 -1479 -89 -1445
rect -147 -1500 -89 -1479
rect -29 1479 29 1500
rect -29 1445 -17 1479
rect 17 1445 29 1479
rect -29 1411 29 1445
rect -29 1377 -17 1411
rect 17 1377 29 1411
rect -29 1343 29 1377
rect -29 1309 -17 1343
rect 17 1309 29 1343
rect -29 1275 29 1309
rect -29 1241 -17 1275
rect 17 1241 29 1275
rect -29 1207 29 1241
rect -29 1173 -17 1207
rect 17 1173 29 1207
rect -29 1139 29 1173
rect -29 1105 -17 1139
rect 17 1105 29 1139
rect -29 1071 29 1105
rect -29 1037 -17 1071
rect 17 1037 29 1071
rect -29 1003 29 1037
rect -29 969 -17 1003
rect 17 969 29 1003
rect -29 935 29 969
rect -29 901 -17 935
rect 17 901 29 935
rect -29 867 29 901
rect -29 833 -17 867
rect 17 833 29 867
rect -29 799 29 833
rect -29 765 -17 799
rect 17 765 29 799
rect -29 731 29 765
rect -29 697 -17 731
rect 17 697 29 731
rect -29 663 29 697
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -697 29 -663
rect -29 -731 -17 -697
rect 17 -731 29 -697
rect -29 -765 29 -731
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -833 29 -799
rect -29 -867 -17 -833
rect 17 -867 29 -833
rect -29 -901 29 -867
rect -29 -935 -17 -901
rect 17 -935 29 -901
rect -29 -969 29 -935
rect -29 -1003 -17 -969
rect 17 -1003 29 -969
rect -29 -1037 29 -1003
rect -29 -1071 -17 -1037
rect 17 -1071 29 -1037
rect -29 -1105 29 -1071
rect -29 -1139 -17 -1105
rect 17 -1139 29 -1105
rect -29 -1173 29 -1139
rect -29 -1207 -17 -1173
rect 17 -1207 29 -1173
rect -29 -1241 29 -1207
rect -29 -1275 -17 -1241
rect 17 -1275 29 -1241
rect -29 -1309 29 -1275
rect -29 -1343 -17 -1309
rect 17 -1343 29 -1309
rect -29 -1377 29 -1343
rect -29 -1411 -17 -1377
rect 17 -1411 29 -1377
rect -29 -1445 29 -1411
rect -29 -1479 -17 -1445
rect 17 -1479 29 -1445
rect -29 -1500 29 -1479
rect 89 1479 147 1500
rect 89 1445 101 1479
rect 135 1445 147 1479
rect 89 1411 147 1445
rect 89 1377 101 1411
rect 135 1377 147 1411
rect 89 1343 147 1377
rect 89 1309 101 1343
rect 135 1309 147 1343
rect 89 1275 147 1309
rect 89 1241 101 1275
rect 135 1241 147 1275
rect 89 1207 147 1241
rect 89 1173 101 1207
rect 135 1173 147 1207
rect 89 1139 147 1173
rect 89 1105 101 1139
rect 135 1105 147 1139
rect 89 1071 147 1105
rect 89 1037 101 1071
rect 135 1037 147 1071
rect 89 1003 147 1037
rect 89 969 101 1003
rect 135 969 147 1003
rect 89 935 147 969
rect 89 901 101 935
rect 135 901 147 935
rect 89 867 147 901
rect 89 833 101 867
rect 135 833 147 867
rect 89 799 147 833
rect 89 765 101 799
rect 135 765 147 799
rect 89 731 147 765
rect 89 697 101 731
rect 135 697 147 731
rect 89 663 147 697
rect 89 629 101 663
rect 135 629 147 663
rect 89 595 147 629
rect 89 561 101 595
rect 135 561 147 595
rect 89 527 147 561
rect 89 493 101 527
rect 135 493 147 527
rect 89 459 147 493
rect 89 425 101 459
rect 135 425 147 459
rect 89 391 147 425
rect 89 357 101 391
rect 135 357 147 391
rect 89 323 147 357
rect 89 289 101 323
rect 135 289 147 323
rect 89 255 147 289
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -289 147 -255
rect 89 -323 101 -289
rect 135 -323 147 -289
rect 89 -357 147 -323
rect 89 -391 101 -357
rect 135 -391 147 -357
rect 89 -425 147 -391
rect 89 -459 101 -425
rect 135 -459 147 -425
rect 89 -493 147 -459
rect 89 -527 101 -493
rect 135 -527 147 -493
rect 89 -561 147 -527
rect 89 -595 101 -561
rect 135 -595 147 -561
rect 89 -629 147 -595
rect 89 -663 101 -629
rect 135 -663 147 -629
rect 89 -697 147 -663
rect 89 -731 101 -697
rect 135 -731 147 -697
rect 89 -765 147 -731
rect 89 -799 101 -765
rect 135 -799 147 -765
rect 89 -833 147 -799
rect 89 -867 101 -833
rect 135 -867 147 -833
rect 89 -901 147 -867
rect 89 -935 101 -901
rect 135 -935 147 -901
rect 89 -969 147 -935
rect 89 -1003 101 -969
rect 135 -1003 147 -969
rect 89 -1037 147 -1003
rect 89 -1071 101 -1037
rect 135 -1071 147 -1037
rect 89 -1105 147 -1071
rect 89 -1139 101 -1105
rect 135 -1139 147 -1105
rect 89 -1173 147 -1139
rect 89 -1207 101 -1173
rect 135 -1207 147 -1173
rect 89 -1241 147 -1207
rect 89 -1275 101 -1241
rect 135 -1275 147 -1241
rect 89 -1309 147 -1275
rect 89 -1343 101 -1309
rect 135 -1343 147 -1309
rect 89 -1377 147 -1343
rect 89 -1411 101 -1377
rect 135 -1411 147 -1377
rect 89 -1445 147 -1411
rect 89 -1479 101 -1445
rect 135 -1479 147 -1445
rect 89 -1500 147 -1479
rect 207 1479 265 1500
rect 207 1445 219 1479
rect 253 1445 265 1479
rect 207 1411 265 1445
rect 207 1377 219 1411
rect 253 1377 265 1411
rect 207 1343 265 1377
rect 207 1309 219 1343
rect 253 1309 265 1343
rect 207 1275 265 1309
rect 207 1241 219 1275
rect 253 1241 265 1275
rect 207 1207 265 1241
rect 207 1173 219 1207
rect 253 1173 265 1207
rect 207 1139 265 1173
rect 207 1105 219 1139
rect 253 1105 265 1139
rect 207 1071 265 1105
rect 207 1037 219 1071
rect 253 1037 265 1071
rect 207 1003 265 1037
rect 207 969 219 1003
rect 253 969 265 1003
rect 207 935 265 969
rect 207 901 219 935
rect 253 901 265 935
rect 207 867 265 901
rect 207 833 219 867
rect 253 833 265 867
rect 207 799 265 833
rect 207 765 219 799
rect 253 765 265 799
rect 207 731 265 765
rect 207 697 219 731
rect 253 697 265 731
rect 207 663 265 697
rect 207 629 219 663
rect 253 629 265 663
rect 207 595 265 629
rect 207 561 219 595
rect 253 561 265 595
rect 207 527 265 561
rect 207 493 219 527
rect 253 493 265 527
rect 207 459 265 493
rect 207 425 219 459
rect 253 425 265 459
rect 207 391 265 425
rect 207 357 219 391
rect 253 357 265 391
rect 207 323 265 357
rect 207 289 219 323
rect 253 289 265 323
rect 207 255 265 289
rect 207 221 219 255
rect 253 221 265 255
rect 207 187 265 221
rect 207 153 219 187
rect 253 153 265 187
rect 207 119 265 153
rect 207 85 219 119
rect 253 85 265 119
rect 207 51 265 85
rect 207 17 219 51
rect 253 17 265 51
rect 207 -17 265 17
rect 207 -51 219 -17
rect 253 -51 265 -17
rect 207 -85 265 -51
rect 207 -119 219 -85
rect 253 -119 265 -85
rect 207 -153 265 -119
rect 207 -187 219 -153
rect 253 -187 265 -153
rect 207 -221 265 -187
rect 207 -255 219 -221
rect 253 -255 265 -221
rect 207 -289 265 -255
rect 207 -323 219 -289
rect 253 -323 265 -289
rect 207 -357 265 -323
rect 207 -391 219 -357
rect 253 -391 265 -357
rect 207 -425 265 -391
rect 207 -459 219 -425
rect 253 -459 265 -425
rect 207 -493 265 -459
rect 207 -527 219 -493
rect 253 -527 265 -493
rect 207 -561 265 -527
rect 207 -595 219 -561
rect 253 -595 265 -561
rect 207 -629 265 -595
rect 207 -663 219 -629
rect 253 -663 265 -629
rect 207 -697 265 -663
rect 207 -731 219 -697
rect 253 -731 265 -697
rect 207 -765 265 -731
rect 207 -799 219 -765
rect 253 -799 265 -765
rect 207 -833 265 -799
rect 207 -867 219 -833
rect 253 -867 265 -833
rect 207 -901 265 -867
rect 207 -935 219 -901
rect 253 -935 265 -901
rect 207 -969 265 -935
rect 207 -1003 219 -969
rect 253 -1003 265 -969
rect 207 -1037 265 -1003
rect 207 -1071 219 -1037
rect 253 -1071 265 -1037
rect 207 -1105 265 -1071
rect 207 -1139 219 -1105
rect 253 -1139 265 -1105
rect 207 -1173 265 -1139
rect 207 -1207 219 -1173
rect 253 -1207 265 -1173
rect 207 -1241 265 -1207
rect 207 -1275 219 -1241
rect 253 -1275 265 -1241
rect 207 -1309 265 -1275
rect 207 -1343 219 -1309
rect 253 -1343 265 -1309
rect 207 -1377 265 -1343
rect 207 -1411 219 -1377
rect 253 -1411 265 -1377
rect 207 -1445 265 -1411
rect 207 -1479 219 -1445
rect 253 -1479 265 -1445
rect 207 -1500 265 -1479
<< pdiffc >>
rect -253 1445 -219 1479
rect -253 1377 -219 1411
rect -253 1309 -219 1343
rect -253 1241 -219 1275
rect -253 1173 -219 1207
rect -253 1105 -219 1139
rect -253 1037 -219 1071
rect -253 969 -219 1003
rect -253 901 -219 935
rect -253 833 -219 867
rect -253 765 -219 799
rect -253 697 -219 731
rect -253 629 -219 663
rect -253 561 -219 595
rect -253 493 -219 527
rect -253 425 -219 459
rect -253 357 -219 391
rect -253 289 -219 323
rect -253 221 -219 255
rect -253 153 -219 187
rect -253 85 -219 119
rect -253 17 -219 51
rect -253 -51 -219 -17
rect -253 -119 -219 -85
rect -253 -187 -219 -153
rect -253 -255 -219 -221
rect -253 -323 -219 -289
rect -253 -391 -219 -357
rect -253 -459 -219 -425
rect -253 -527 -219 -493
rect -253 -595 -219 -561
rect -253 -663 -219 -629
rect -253 -731 -219 -697
rect -253 -799 -219 -765
rect -253 -867 -219 -833
rect -253 -935 -219 -901
rect -253 -1003 -219 -969
rect -253 -1071 -219 -1037
rect -253 -1139 -219 -1105
rect -253 -1207 -219 -1173
rect -253 -1275 -219 -1241
rect -253 -1343 -219 -1309
rect -253 -1411 -219 -1377
rect -253 -1479 -219 -1445
rect -135 1445 -101 1479
rect -135 1377 -101 1411
rect -135 1309 -101 1343
rect -135 1241 -101 1275
rect -135 1173 -101 1207
rect -135 1105 -101 1139
rect -135 1037 -101 1071
rect -135 969 -101 1003
rect -135 901 -101 935
rect -135 833 -101 867
rect -135 765 -101 799
rect -135 697 -101 731
rect -135 629 -101 663
rect -135 561 -101 595
rect -135 493 -101 527
rect -135 425 -101 459
rect -135 357 -101 391
rect -135 289 -101 323
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -135 -323 -101 -289
rect -135 -391 -101 -357
rect -135 -459 -101 -425
rect -135 -527 -101 -493
rect -135 -595 -101 -561
rect -135 -663 -101 -629
rect -135 -731 -101 -697
rect -135 -799 -101 -765
rect -135 -867 -101 -833
rect -135 -935 -101 -901
rect -135 -1003 -101 -969
rect -135 -1071 -101 -1037
rect -135 -1139 -101 -1105
rect -135 -1207 -101 -1173
rect -135 -1275 -101 -1241
rect -135 -1343 -101 -1309
rect -135 -1411 -101 -1377
rect -135 -1479 -101 -1445
rect -17 1445 17 1479
rect -17 1377 17 1411
rect -17 1309 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1139
rect -17 1037 17 1071
rect -17 969 17 1003
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1003 17 -969
rect -17 -1071 17 -1037
rect -17 -1139 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1309
rect -17 -1411 17 -1377
rect -17 -1479 17 -1445
rect 101 1445 135 1479
rect 101 1377 135 1411
rect 101 1309 135 1343
rect 101 1241 135 1275
rect 101 1173 135 1207
rect 101 1105 135 1139
rect 101 1037 135 1071
rect 101 969 135 1003
rect 101 901 135 935
rect 101 833 135 867
rect 101 765 135 799
rect 101 697 135 731
rect 101 629 135 663
rect 101 561 135 595
rect 101 493 135 527
rect 101 425 135 459
rect 101 357 135 391
rect 101 289 135 323
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
rect 101 -323 135 -289
rect 101 -391 135 -357
rect 101 -459 135 -425
rect 101 -527 135 -493
rect 101 -595 135 -561
rect 101 -663 135 -629
rect 101 -731 135 -697
rect 101 -799 135 -765
rect 101 -867 135 -833
rect 101 -935 135 -901
rect 101 -1003 135 -969
rect 101 -1071 135 -1037
rect 101 -1139 135 -1105
rect 101 -1207 135 -1173
rect 101 -1275 135 -1241
rect 101 -1343 135 -1309
rect 101 -1411 135 -1377
rect 101 -1479 135 -1445
rect 219 1445 253 1479
rect 219 1377 253 1411
rect 219 1309 253 1343
rect 219 1241 253 1275
rect 219 1173 253 1207
rect 219 1105 253 1139
rect 219 1037 253 1071
rect 219 969 253 1003
rect 219 901 253 935
rect 219 833 253 867
rect 219 765 253 799
rect 219 697 253 731
rect 219 629 253 663
rect 219 561 253 595
rect 219 493 253 527
rect 219 425 253 459
rect 219 357 253 391
rect 219 289 253 323
rect 219 221 253 255
rect 219 153 253 187
rect 219 85 253 119
rect 219 17 253 51
rect 219 -51 253 -17
rect 219 -119 253 -85
rect 219 -187 253 -153
rect 219 -255 253 -221
rect 219 -323 253 -289
rect 219 -391 253 -357
rect 219 -459 253 -425
rect 219 -527 253 -493
rect 219 -595 253 -561
rect 219 -663 253 -629
rect 219 -731 253 -697
rect 219 -799 253 -765
rect 219 -867 253 -833
rect 219 -935 253 -901
rect 219 -1003 253 -969
rect 219 -1071 253 -1037
rect 219 -1139 253 -1105
rect 219 -1207 253 -1173
rect 219 -1275 253 -1241
rect 219 -1343 253 -1309
rect 219 -1411 253 -1377
rect 219 -1479 253 -1445
<< nsubdiff >>
rect -367 1649 -255 1683
rect -221 1649 -187 1683
rect -153 1649 -119 1683
rect -85 1649 -51 1683
rect -17 1649 17 1683
rect 51 1649 85 1683
rect 119 1649 153 1683
rect 187 1649 221 1683
rect 255 1649 367 1683
rect -367 1581 -333 1649
rect -367 1513 -333 1547
rect 333 1581 367 1649
rect 333 1513 367 1547
rect -367 1445 -333 1479
rect -367 1377 -333 1411
rect -367 1309 -333 1343
rect -367 1241 -333 1275
rect -367 1173 -333 1207
rect -367 1105 -333 1139
rect -367 1037 -333 1071
rect -367 969 -333 1003
rect -367 901 -333 935
rect -367 833 -333 867
rect -367 765 -333 799
rect -367 697 -333 731
rect -367 629 -333 663
rect -367 561 -333 595
rect -367 493 -333 527
rect -367 425 -333 459
rect -367 357 -333 391
rect -367 289 -333 323
rect -367 221 -333 255
rect -367 153 -333 187
rect -367 85 -333 119
rect -367 17 -333 51
rect -367 -51 -333 -17
rect -367 -119 -333 -85
rect -367 -187 -333 -153
rect -367 -255 -333 -221
rect -367 -323 -333 -289
rect -367 -391 -333 -357
rect -367 -459 -333 -425
rect -367 -527 -333 -493
rect -367 -595 -333 -561
rect -367 -663 -333 -629
rect -367 -731 -333 -697
rect -367 -799 -333 -765
rect -367 -867 -333 -833
rect -367 -935 -333 -901
rect -367 -1003 -333 -969
rect -367 -1071 -333 -1037
rect -367 -1139 -333 -1105
rect -367 -1207 -333 -1173
rect -367 -1275 -333 -1241
rect -367 -1343 -333 -1309
rect -367 -1411 -333 -1377
rect -367 -1479 -333 -1445
rect 333 1445 367 1479
rect 333 1377 367 1411
rect 333 1309 367 1343
rect 333 1241 367 1275
rect 333 1173 367 1207
rect 333 1105 367 1139
rect 333 1037 367 1071
rect 333 969 367 1003
rect 333 901 367 935
rect 333 833 367 867
rect 333 765 367 799
rect 333 697 367 731
rect 333 629 367 663
rect 333 561 367 595
rect 333 493 367 527
rect 333 425 367 459
rect 333 357 367 391
rect 333 289 367 323
rect 333 221 367 255
rect 333 153 367 187
rect 333 85 367 119
rect 333 17 367 51
rect 333 -51 367 -17
rect 333 -119 367 -85
rect 333 -187 367 -153
rect 333 -255 367 -221
rect 333 -323 367 -289
rect 333 -391 367 -357
rect 333 -459 367 -425
rect 333 -527 367 -493
rect 333 -595 367 -561
rect 333 -663 367 -629
rect 333 -731 367 -697
rect 333 -799 367 -765
rect 333 -867 367 -833
rect 333 -935 367 -901
rect 333 -1003 367 -969
rect 333 -1071 367 -1037
rect 333 -1139 367 -1105
rect 333 -1207 367 -1173
rect 333 -1275 367 -1241
rect 333 -1343 367 -1309
rect 333 -1411 367 -1377
rect 333 -1479 367 -1445
rect -367 -1547 -333 -1513
rect -367 -1649 -333 -1581
rect 333 -1547 367 -1513
rect 333 -1649 367 -1581
rect -367 -1683 -255 -1649
rect -221 -1683 -187 -1649
rect -153 -1683 -119 -1649
rect -85 -1683 -51 -1649
rect -17 -1683 17 -1649
rect 51 -1683 85 -1649
rect 119 -1683 153 -1649
rect 187 -1683 221 -1649
rect 255 -1683 367 -1649
<< nsubdiffcont >>
rect -255 1649 -221 1683
rect -187 1649 -153 1683
rect -119 1649 -85 1683
rect -51 1649 -17 1683
rect 17 1649 51 1683
rect 85 1649 119 1683
rect 153 1649 187 1683
rect 221 1649 255 1683
rect -367 1547 -333 1581
rect 333 1547 367 1581
rect -367 1479 -333 1513
rect -367 1411 -333 1445
rect -367 1343 -333 1377
rect -367 1275 -333 1309
rect -367 1207 -333 1241
rect -367 1139 -333 1173
rect -367 1071 -333 1105
rect -367 1003 -333 1037
rect -367 935 -333 969
rect -367 867 -333 901
rect -367 799 -333 833
rect -367 731 -333 765
rect -367 663 -333 697
rect -367 595 -333 629
rect -367 527 -333 561
rect -367 459 -333 493
rect -367 391 -333 425
rect -367 323 -333 357
rect -367 255 -333 289
rect -367 187 -333 221
rect -367 119 -333 153
rect -367 51 -333 85
rect -367 -17 -333 17
rect -367 -85 -333 -51
rect -367 -153 -333 -119
rect -367 -221 -333 -187
rect -367 -289 -333 -255
rect -367 -357 -333 -323
rect -367 -425 -333 -391
rect -367 -493 -333 -459
rect -367 -561 -333 -527
rect -367 -629 -333 -595
rect -367 -697 -333 -663
rect -367 -765 -333 -731
rect -367 -833 -333 -799
rect -367 -901 -333 -867
rect -367 -969 -333 -935
rect -367 -1037 -333 -1003
rect -367 -1105 -333 -1071
rect -367 -1173 -333 -1139
rect -367 -1241 -333 -1207
rect -367 -1309 -333 -1275
rect -367 -1377 -333 -1343
rect -367 -1445 -333 -1411
rect -367 -1513 -333 -1479
rect 333 1479 367 1513
rect 333 1411 367 1445
rect 333 1343 367 1377
rect 333 1275 367 1309
rect 333 1207 367 1241
rect 333 1139 367 1173
rect 333 1071 367 1105
rect 333 1003 367 1037
rect 333 935 367 969
rect 333 867 367 901
rect 333 799 367 833
rect 333 731 367 765
rect 333 663 367 697
rect 333 595 367 629
rect 333 527 367 561
rect 333 459 367 493
rect 333 391 367 425
rect 333 323 367 357
rect 333 255 367 289
rect 333 187 367 221
rect 333 119 367 153
rect 333 51 367 85
rect 333 -17 367 17
rect 333 -85 367 -51
rect 333 -153 367 -119
rect 333 -221 367 -187
rect 333 -289 367 -255
rect 333 -357 367 -323
rect 333 -425 367 -391
rect 333 -493 367 -459
rect 333 -561 367 -527
rect 333 -629 367 -595
rect 333 -697 367 -663
rect 333 -765 367 -731
rect 333 -833 367 -799
rect 333 -901 367 -867
rect 333 -969 367 -935
rect 333 -1037 367 -1003
rect 333 -1105 367 -1071
rect 333 -1173 367 -1139
rect 333 -1241 367 -1207
rect 333 -1309 367 -1275
rect 333 -1377 367 -1343
rect 333 -1445 367 -1411
rect 333 -1513 367 -1479
rect -367 -1581 -333 -1547
rect 333 -1581 367 -1547
rect -255 -1683 -221 -1649
rect -187 -1683 -153 -1649
rect -119 -1683 -85 -1649
rect -51 -1683 -17 -1649
rect 17 -1683 51 -1649
rect 85 -1683 119 -1649
rect 153 -1683 187 -1649
rect 221 -1683 255 -1649
<< poly >>
rect -210 1581 -144 1597
rect -210 1547 -194 1581
rect -160 1547 -144 1581
rect -210 1531 -144 1547
rect -92 1581 -26 1597
rect -92 1547 -76 1581
rect -42 1547 -26 1581
rect -92 1531 -26 1547
rect 26 1581 92 1597
rect 26 1547 42 1581
rect 76 1547 92 1581
rect 26 1531 92 1547
rect 144 1581 210 1597
rect 144 1547 160 1581
rect 194 1547 210 1581
rect 144 1531 210 1547
rect -207 1500 -147 1531
rect -89 1500 -29 1531
rect 29 1500 89 1531
rect 147 1500 207 1531
rect -207 -1531 -147 -1500
rect -89 -1531 -29 -1500
rect 29 -1531 89 -1500
rect 147 -1531 207 -1500
rect -210 -1547 -144 -1531
rect -210 -1581 -194 -1547
rect -160 -1581 -144 -1547
rect -210 -1597 -144 -1581
rect -92 -1547 -26 -1531
rect -92 -1581 -76 -1547
rect -42 -1581 -26 -1547
rect -92 -1597 -26 -1581
rect 26 -1547 92 -1531
rect 26 -1581 42 -1547
rect 76 -1581 92 -1547
rect 26 -1597 92 -1581
rect 144 -1547 210 -1531
rect 144 -1581 160 -1547
rect 194 -1581 210 -1547
rect 144 -1597 210 -1581
<< polycont >>
rect -194 1547 -160 1581
rect -76 1547 -42 1581
rect 42 1547 76 1581
rect 160 1547 194 1581
rect -194 -1581 -160 -1547
rect -76 -1581 -42 -1547
rect 42 -1581 76 -1547
rect 160 -1581 194 -1547
<< locali >>
rect -367 1649 -255 1683
rect -221 1649 -187 1683
rect -153 1649 -119 1683
rect -85 1649 -51 1683
rect -17 1649 17 1683
rect 51 1649 85 1683
rect 119 1649 153 1683
rect 187 1649 221 1683
rect 255 1649 367 1683
rect -367 1581 -333 1649
rect 333 1581 367 1649
rect -210 1547 -194 1581
rect -160 1547 -144 1581
rect -92 1547 -76 1581
rect -42 1547 -26 1581
rect 26 1547 42 1581
rect 76 1547 92 1581
rect 144 1547 160 1581
rect 194 1547 210 1581
rect -367 1513 -333 1547
rect 333 1513 367 1547
rect -367 1445 -333 1479
rect -367 1377 -333 1411
rect -367 1309 -333 1343
rect -367 1241 -333 1275
rect -367 1173 -333 1207
rect -367 1105 -333 1139
rect -367 1037 -333 1071
rect -367 969 -333 1003
rect -367 901 -333 935
rect -367 833 -333 867
rect -367 765 -333 799
rect -367 697 -333 731
rect -367 629 -333 663
rect -367 561 -333 595
rect -367 493 -333 527
rect -367 425 -333 459
rect -367 357 -333 391
rect -367 289 -333 323
rect -367 221 -333 255
rect -367 153 -333 187
rect -367 85 -333 119
rect -367 17 -333 51
rect -367 -51 -333 -17
rect -367 -119 -333 -85
rect -367 -187 -333 -153
rect -367 -255 -333 -221
rect -367 -323 -333 -289
rect -367 -391 -333 -357
rect -367 -459 -333 -425
rect -367 -527 -333 -493
rect -367 -595 -333 -561
rect -367 -663 -333 -629
rect -367 -731 -333 -697
rect -367 -799 -333 -765
rect -367 -867 -333 -833
rect -367 -935 -333 -901
rect -367 -1003 -333 -969
rect -367 -1071 -333 -1037
rect -367 -1139 -333 -1105
rect -367 -1207 -333 -1173
rect -367 -1275 -333 -1241
rect -367 -1343 -333 -1309
rect -367 -1411 -333 -1377
rect -367 -1479 -333 -1445
rect -253 1479 -219 1504
rect -253 1411 -219 1423
rect -253 1343 -219 1351
rect -253 1275 -219 1279
rect -253 1169 -219 1173
rect -253 1097 -219 1105
rect -253 1025 -219 1037
rect -253 953 -219 969
rect -253 881 -219 901
rect -253 809 -219 833
rect -253 737 -219 765
rect -253 665 -219 697
rect -253 595 -219 629
rect -253 527 -219 559
rect -253 459 -219 487
rect -253 391 -219 415
rect -253 323 -219 343
rect -253 255 -219 271
rect -253 187 -219 199
rect -253 119 -219 127
rect -253 51 -219 55
rect -253 -55 -219 -51
rect -253 -127 -219 -119
rect -253 -199 -219 -187
rect -253 -271 -219 -255
rect -253 -343 -219 -323
rect -253 -415 -219 -391
rect -253 -487 -219 -459
rect -253 -559 -219 -527
rect -253 -629 -219 -595
rect -253 -697 -219 -665
rect -253 -765 -219 -737
rect -253 -833 -219 -809
rect -253 -901 -219 -881
rect -253 -969 -219 -953
rect -253 -1037 -219 -1025
rect -253 -1105 -219 -1097
rect -253 -1173 -219 -1169
rect -253 -1279 -219 -1275
rect -253 -1351 -219 -1343
rect -253 -1423 -219 -1411
rect -253 -1504 -219 -1479
rect -135 1479 -101 1504
rect -135 1411 -101 1423
rect -135 1343 -101 1351
rect -135 1275 -101 1279
rect -135 1169 -101 1173
rect -135 1097 -101 1105
rect -135 1025 -101 1037
rect -135 953 -101 969
rect -135 881 -101 901
rect -135 809 -101 833
rect -135 737 -101 765
rect -135 665 -101 697
rect -135 595 -101 629
rect -135 527 -101 559
rect -135 459 -101 487
rect -135 391 -101 415
rect -135 323 -101 343
rect -135 255 -101 271
rect -135 187 -101 199
rect -135 119 -101 127
rect -135 51 -101 55
rect -135 -55 -101 -51
rect -135 -127 -101 -119
rect -135 -199 -101 -187
rect -135 -271 -101 -255
rect -135 -343 -101 -323
rect -135 -415 -101 -391
rect -135 -487 -101 -459
rect -135 -559 -101 -527
rect -135 -629 -101 -595
rect -135 -697 -101 -665
rect -135 -765 -101 -737
rect -135 -833 -101 -809
rect -135 -901 -101 -881
rect -135 -969 -101 -953
rect -135 -1037 -101 -1025
rect -135 -1105 -101 -1097
rect -135 -1173 -101 -1169
rect -135 -1279 -101 -1275
rect -135 -1351 -101 -1343
rect -135 -1423 -101 -1411
rect -135 -1504 -101 -1479
rect -17 1479 17 1504
rect -17 1411 17 1423
rect -17 1343 17 1351
rect -17 1275 17 1279
rect -17 1169 17 1173
rect -17 1097 17 1105
rect -17 1025 17 1037
rect -17 953 17 969
rect -17 881 17 901
rect -17 809 17 833
rect -17 737 17 765
rect -17 665 17 697
rect -17 595 17 629
rect -17 527 17 559
rect -17 459 17 487
rect -17 391 17 415
rect -17 323 17 343
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -343 17 -323
rect -17 -415 17 -391
rect -17 -487 17 -459
rect -17 -559 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -665
rect -17 -765 17 -737
rect -17 -833 17 -809
rect -17 -901 17 -881
rect -17 -969 17 -953
rect -17 -1037 17 -1025
rect -17 -1105 17 -1097
rect -17 -1173 17 -1169
rect -17 -1279 17 -1275
rect -17 -1351 17 -1343
rect -17 -1423 17 -1411
rect -17 -1504 17 -1479
rect 101 1479 135 1504
rect 101 1411 135 1423
rect 101 1343 135 1351
rect 101 1275 135 1279
rect 101 1169 135 1173
rect 101 1097 135 1105
rect 101 1025 135 1037
rect 101 953 135 969
rect 101 881 135 901
rect 101 809 135 833
rect 101 737 135 765
rect 101 665 135 697
rect 101 595 135 629
rect 101 527 135 559
rect 101 459 135 487
rect 101 391 135 415
rect 101 323 135 343
rect 101 255 135 271
rect 101 187 135 199
rect 101 119 135 127
rect 101 51 135 55
rect 101 -55 135 -51
rect 101 -127 135 -119
rect 101 -199 135 -187
rect 101 -271 135 -255
rect 101 -343 135 -323
rect 101 -415 135 -391
rect 101 -487 135 -459
rect 101 -559 135 -527
rect 101 -629 135 -595
rect 101 -697 135 -665
rect 101 -765 135 -737
rect 101 -833 135 -809
rect 101 -901 135 -881
rect 101 -969 135 -953
rect 101 -1037 135 -1025
rect 101 -1105 135 -1097
rect 101 -1173 135 -1169
rect 101 -1279 135 -1275
rect 101 -1351 135 -1343
rect 101 -1423 135 -1411
rect 101 -1504 135 -1479
rect 219 1479 253 1504
rect 219 1411 253 1423
rect 219 1343 253 1351
rect 219 1275 253 1279
rect 219 1169 253 1173
rect 219 1097 253 1105
rect 219 1025 253 1037
rect 219 953 253 969
rect 219 881 253 901
rect 219 809 253 833
rect 219 737 253 765
rect 219 665 253 697
rect 219 595 253 629
rect 219 527 253 559
rect 219 459 253 487
rect 219 391 253 415
rect 219 323 253 343
rect 219 255 253 271
rect 219 187 253 199
rect 219 119 253 127
rect 219 51 253 55
rect 219 -55 253 -51
rect 219 -127 253 -119
rect 219 -199 253 -187
rect 219 -271 253 -255
rect 219 -343 253 -323
rect 219 -415 253 -391
rect 219 -487 253 -459
rect 219 -559 253 -527
rect 219 -629 253 -595
rect 219 -697 253 -665
rect 219 -765 253 -737
rect 219 -833 253 -809
rect 219 -901 253 -881
rect 219 -969 253 -953
rect 219 -1037 253 -1025
rect 219 -1105 253 -1097
rect 219 -1173 253 -1169
rect 219 -1279 253 -1275
rect 219 -1351 253 -1343
rect 219 -1423 253 -1411
rect 219 -1504 253 -1479
rect 333 1445 367 1479
rect 333 1377 367 1411
rect 333 1309 367 1343
rect 333 1241 367 1275
rect 333 1173 367 1207
rect 333 1105 367 1139
rect 333 1037 367 1071
rect 333 969 367 1003
rect 333 901 367 935
rect 333 833 367 867
rect 333 765 367 799
rect 333 697 367 731
rect 333 629 367 663
rect 333 561 367 595
rect 333 493 367 527
rect 333 425 367 459
rect 333 357 367 391
rect 333 289 367 323
rect 333 221 367 255
rect 333 153 367 187
rect 333 85 367 119
rect 333 17 367 51
rect 333 -51 367 -17
rect 333 -119 367 -85
rect 333 -187 367 -153
rect 333 -255 367 -221
rect 333 -323 367 -289
rect 333 -391 367 -357
rect 333 -459 367 -425
rect 333 -527 367 -493
rect 333 -595 367 -561
rect 333 -663 367 -629
rect 333 -731 367 -697
rect 333 -799 367 -765
rect 333 -867 367 -833
rect 333 -935 367 -901
rect 333 -1003 367 -969
rect 333 -1071 367 -1037
rect 333 -1139 367 -1105
rect 333 -1207 367 -1173
rect 333 -1275 367 -1241
rect 333 -1343 367 -1309
rect 333 -1411 367 -1377
rect 333 -1479 367 -1445
rect -367 -1547 -333 -1513
rect 333 -1547 367 -1513
rect -210 -1581 -194 -1547
rect -160 -1581 -144 -1547
rect -92 -1581 -76 -1547
rect -42 -1581 -26 -1547
rect 26 -1581 42 -1547
rect 76 -1581 92 -1547
rect 144 -1581 160 -1547
rect 194 -1581 210 -1547
rect -367 -1649 -333 -1581
rect 333 -1649 367 -1581
rect -367 -1683 -255 -1649
rect -221 -1683 -187 -1649
rect -153 -1683 -119 -1649
rect -85 -1683 -51 -1649
rect -17 -1683 17 -1649
rect 51 -1683 85 -1649
rect 119 -1683 153 -1649
rect 187 -1683 221 -1649
rect 255 -1683 367 -1649
<< viali >>
rect -194 1547 -160 1581
rect -76 1547 -42 1581
rect 42 1547 76 1581
rect 160 1547 194 1581
rect -253 1445 -219 1457
rect -253 1423 -219 1445
rect -253 1377 -219 1385
rect -253 1351 -219 1377
rect -253 1309 -219 1313
rect -253 1279 -219 1309
rect -253 1207 -219 1241
rect -253 1139 -219 1169
rect -253 1135 -219 1139
rect -253 1071 -219 1097
rect -253 1063 -219 1071
rect -253 1003 -219 1025
rect -253 991 -219 1003
rect -253 935 -219 953
rect -253 919 -219 935
rect -253 867 -219 881
rect -253 847 -219 867
rect -253 799 -219 809
rect -253 775 -219 799
rect -253 731 -219 737
rect -253 703 -219 731
rect -253 663 -219 665
rect -253 631 -219 663
rect -253 561 -219 593
rect -253 559 -219 561
rect -253 493 -219 521
rect -253 487 -219 493
rect -253 425 -219 449
rect -253 415 -219 425
rect -253 357 -219 377
rect -253 343 -219 357
rect -253 289 -219 305
rect -253 271 -219 289
rect -253 221 -219 233
rect -253 199 -219 221
rect -253 153 -219 161
rect -253 127 -219 153
rect -253 85 -219 89
rect -253 55 -219 85
rect -253 -17 -219 17
rect -253 -85 -219 -55
rect -253 -89 -219 -85
rect -253 -153 -219 -127
rect -253 -161 -219 -153
rect -253 -221 -219 -199
rect -253 -233 -219 -221
rect -253 -289 -219 -271
rect -253 -305 -219 -289
rect -253 -357 -219 -343
rect -253 -377 -219 -357
rect -253 -425 -219 -415
rect -253 -449 -219 -425
rect -253 -493 -219 -487
rect -253 -521 -219 -493
rect -253 -561 -219 -559
rect -253 -593 -219 -561
rect -253 -663 -219 -631
rect -253 -665 -219 -663
rect -253 -731 -219 -703
rect -253 -737 -219 -731
rect -253 -799 -219 -775
rect -253 -809 -219 -799
rect -253 -867 -219 -847
rect -253 -881 -219 -867
rect -253 -935 -219 -919
rect -253 -953 -219 -935
rect -253 -1003 -219 -991
rect -253 -1025 -219 -1003
rect -253 -1071 -219 -1063
rect -253 -1097 -219 -1071
rect -253 -1139 -219 -1135
rect -253 -1169 -219 -1139
rect -253 -1241 -219 -1207
rect -253 -1309 -219 -1279
rect -253 -1313 -219 -1309
rect -253 -1377 -219 -1351
rect -253 -1385 -219 -1377
rect -253 -1445 -219 -1423
rect -253 -1457 -219 -1445
rect -135 1445 -101 1457
rect -135 1423 -101 1445
rect -135 1377 -101 1385
rect -135 1351 -101 1377
rect -135 1309 -101 1313
rect -135 1279 -101 1309
rect -135 1207 -101 1241
rect -135 1139 -101 1169
rect -135 1135 -101 1139
rect -135 1071 -101 1097
rect -135 1063 -101 1071
rect -135 1003 -101 1025
rect -135 991 -101 1003
rect -135 935 -101 953
rect -135 919 -101 935
rect -135 867 -101 881
rect -135 847 -101 867
rect -135 799 -101 809
rect -135 775 -101 799
rect -135 731 -101 737
rect -135 703 -101 731
rect -135 663 -101 665
rect -135 631 -101 663
rect -135 561 -101 593
rect -135 559 -101 561
rect -135 493 -101 521
rect -135 487 -101 493
rect -135 425 -101 449
rect -135 415 -101 425
rect -135 357 -101 377
rect -135 343 -101 357
rect -135 289 -101 305
rect -135 271 -101 289
rect -135 221 -101 233
rect -135 199 -101 221
rect -135 153 -101 161
rect -135 127 -101 153
rect -135 85 -101 89
rect -135 55 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -55
rect -135 -89 -101 -85
rect -135 -153 -101 -127
rect -135 -161 -101 -153
rect -135 -221 -101 -199
rect -135 -233 -101 -221
rect -135 -289 -101 -271
rect -135 -305 -101 -289
rect -135 -357 -101 -343
rect -135 -377 -101 -357
rect -135 -425 -101 -415
rect -135 -449 -101 -425
rect -135 -493 -101 -487
rect -135 -521 -101 -493
rect -135 -561 -101 -559
rect -135 -593 -101 -561
rect -135 -663 -101 -631
rect -135 -665 -101 -663
rect -135 -731 -101 -703
rect -135 -737 -101 -731
rect -135 -799 -101 -775
rect -135 -809 -101 -799
rect -135 -867 -101 -847
rect -135 -881 -101 -867
rect -135 -935 -101 -919
rect -135 -953 -101 -935
rect -135 -1003 -101 -991
rect -135 -1025 -101 -1003
rect -135 -1071 -101 -1063
rect -135 -1097 -101 -1071
rect -135 -1139 -101 -1135
rect -135 -1169 -101 -1139
rect -135 -1241 -101 -1207
rect -135 -1309 -101 -1279
rect -135 -1313 -101 -1309
rect -135 -1377 -101 -1351
rect -135 -1385 -101 -1377
rect -135 -1445 -101 -1423
rect -135 -1457 -101 -1445
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect 101 1445 135 1457
rect 101 1423 135 1445
rect 101 1377 135 1385
rect 101 1351 135 1377
rect 101 1309 135 1313
rect 101 1279 135 1309
rect 101 1207 135 1241
rect 101 1139 135 1169
rect 101 1135 135 1139
rect 101 1071 135 1097
rect 101 1063 135 1071
rect 101 1003 135 1025
rect 101 991 135 1003
rect 101 935 135 953
rect 101 919 135 935
rect 101 867 135 881
rect 101 847 135 867
rect 101 799 135 809
rect 101 775 135 799
rect 101 731 135 737
rect 101 703 135 731
rect 101 663 135 665
rect 101 631 135 663
rect 101 561 135 593
rect 101 559 135 561
rect 101 493 135 521
rect 101 487 135 493
rect 101 425 135 449
rect 101 415 135 425
rect 101 357 135 377
rect 101 343 135 357
rect 101 289 135 305
rect 101 271 135 289
rect 101 221 135 233
rect 101 199 135 221
rect 101 153 135 161
rect 101 127 135 153
rect 101 85 135 89
rect 101 55 135 85
rect 101 -17 135 17
rect 101 -85 135 -55
rect 101 -89 135 -85
rect 101 -153 135 -127
rect 101 -161 135 -153
rect 101 -221 135 -199
rect 101 -233 135 -221
rect 101 -289 135 -271
rect 101 -305 135 -289
rect 101 -357 135 -343
rect 101 -377 135 -357
rect 101 -425 135 -415
rect 101 -449 135 -425
rect 101 -493 135 -487
rect 101 -521 135 -493
rect 101 -561 135 -559
rect 101 -593 135 -561
rect 101 -663 135 -631
rect 101 -665 135 -663
rect 101 -731 135 -703
rect 101 -737 135 -731
rect 101 -799 135 -775
rect 101 -809 135 -799
rect 101 -867 135 -847
rect 101 -881 135 -867
rect 101 -935 135 -919
rect 101 -953 135 -935
rect 101 -1003 135 -991
rect 101 -1025 135 -1003
rect 101 -1071 135 -1063
rect 101 -1097 135 -1071
rect 101 -1139 135 -1135
rect 101 -1169 135 -1139
rect 101 -1241 135 -1207
rect 101 -1309 135 -1279
rect 101 -1313 135 -1309
rect 101 -1377 135 -1351
rect 101 -1385 135 -1377
rect 101 -1445 135 -1423
rect 101 -1457 135 -1445
rect 219 1445 253 1457
rect 219 1423 253 1445
rect 219 1377 253 1385
rect 219 1351 253 1377
rect 219 1309 253 1313
rect 219 1279 253 1309
rect 219 1207 253 1241
rect 219 1139 253 1169
rect 219 1135 253 1139
rect 219 1071 253 1097
rect 219 1063 253 1071
rect 219 1003 253 1025
rect 219 991 253 1003
rect 219 935 253 953
rect 219 919 253 935
rect 219 867 253 881
rect 219 847 253 867
rect 219 799 253 809
rect 219 775 253 799
rect 219 731 253 737
rect 219 703 253 731
rect 219 663 253 665
rect 219 631 253 663
rect 219 561 253 593
rect 219 559 253 561
rect 219 493 253 521
rect 219 487 253 493
rect 219 425 253 449
rect 219 415 253 425
rect 219 357 253 377
rect 219 343 253 357
rect 219 289 253 305
rect 219 271 253 289
rect 219 221 253 233
rect 219 199 253 221
rect 219 153 253 161
rect 219 127 253 153
rect 219 85 253 89
rect 219 55 253 85
rect 219 -17 253 17
rect 219 -85 253 -55
rect 219 -89 253 -85
rect 219 -153 253 -127
rect 219 -161 253 -153
rect 219 -221 253 -199
rect 219 -233 253 -221
rect 219 -289 253 -271
rect 219 -305 253 -289
rect 219 -357 253 -343
rect 219 -377 253 -357
rect 219 -425 253 -415
rect 219 -449 253 -425
rect 219 -493 253 -487
rect 219 -521 253 -493
rect 219 -561 253 -559
rect 219 -593 253 -561
rect 219 -663 253 -631
rect 219 -665 253 -663
rect 219 -731 253 -703
rect 219 -737 253 -731
rect 219 -799 253 -775
rect 219 -809 253 -799
rect 219 -867 253 -847
rect 219 -881 253 -867
rect 219 -935 253 -919
rect 219 -953 253 -935
rect 219 -1003 253 -991
rect 219 -1025 253 -1003
rect 219 -1071 253 -1063
rect 219 -1097 253 -1071
rect 219 -1139 253 -1135
rect 219 -1169 253 -1139
rect 219 -1241 253 -1207
rect 219 -1309 253 -1279
rect 219 -1313 253 -1309
rect 219 -1377 253 -1351
rect 219 -1385 253 -1377
rect 219 -1445 253 -1423
rect 219 -1457 253 -1445
rect -194 -1581 -160 -1547
rect -76 -1581 -42 -1547
rect 42 -1581 76 -1547
rect 160 -1581 194 -1547
<< metal1 >>
rect -206 1581 -148 1587
rect -206 1547 -194 1581
rect -160 1547 -148 1581
rect -206 1541 -148 1547
rect -88 1581 -30 1587
rect -88 1547 -76 1581
rect -42 1547 -30 1581
rect -88 1541 -30 1547
rect 30 1581 88 1587
rect 30 1547 42 1581
rect 76 1547 88 1581
rect 30 1541 88 1547
rect 148 1581 206 1587
rect 148 1547 160 1581
rect 194 1547 206 1581
rect 148 1541 206 1547
rect -259 1457 -213 1500
rect -259 1423 -253 1457
rect -219 1423 -213 1457
rect -259 1385 -213 1423
rect -259 1351 -253 1385
rect -219 1351 -213 1385
rect -259 1313 -213 1351
rect -259 1279 -253 1313
rect -219 1279 -213 1313
rect -259 1241 -213 1279
rect -259 1207 -253 1241
rect -219 1207 -213 1241
rect -259 1169 -213 1207
rect -259 1135 -253 1169
rect -219 1135 -213 1169
rect -259 1097 -213 1135
rect -259 1063 -253 1097
rect -219 1063 -213 1097
rect -259 1025 -213 1063
rect -259 991 -253 1025
rect -219 991 -213 1025
rect -259 953 -213 991
rect -259 919 -253 953
rect -219 919 -213 953
rect -259 881 -213 919
rect -259 847 -253 881
rect -219 847 -213 881
rect -259 809 -213 847
rect -259 775 -253 809
rect -219 775 -213 809
rect -259 737 -213 775
rect -259 703 -253 737
rect -219 703 -213 737
rect -259 665 -213 703
rect -259 631 -253 665
rect -219 631 -213 665
rect -259 593 -213 631
rect -259 559 -253 593
rect -219 559 -213 593
rect -259 521 -213 559
rect -259 487 -253 521
rect -219 487 -213 521
rect -259 449 -213 487
rect -259 415 -253 449
rect -219 415 -213 449
rect -259 377 -213 415
rect -259 343 -253 377
rect -219 343 -213 377
rect -259 305 -213 343
rect -259 271 -253 305
rect -219 271 -213 305
rect -259 233 -213 271
rect -259 199 -253 233
rect -219 199 -213 233
rect -259 161 -213 199
rect -259 127 -253 161
rect -219 127 -213 161
rect -259 89 -213 127
rect -259 55 -253 89
rect -219 55 -213 89
rect -259 17 -213 55
rect -259 -17 -253 17
rect -219 -17 -213 17
rect -259 -55 -213 -17
rect -259 -89 -253 -55
rect -219 -89 -213 -55
rect -259 -127 -213 -89
rect -259 -161 -253 -127
rect -219 -161 -213 -127
rect -259 -199 -213 -161
rect -259 -233 -253 -199
rect -219 -233 -213 -199
rect -259 -271 -213 -233
rect -259 -305 -253 -271
rect -219 -305 -213 -271
rect -259 -343 -213 -305
rect -259 -377 -253 -343
rect -219 -377 -213 -343
rect -259 -415 -213 -377
rect -259 -449 -253 -415
rect -219 -449 -213 -415
rect -259 -487 -213 -449
rect -259 -521 -253 -487
rect -219 -521 -213 -487
rect -259 -559 -213 -521
rect -259 -593 -253 -559
rect -219 -593 -213 -559
rect -259 -631 -213 -593
rect -259 -665 -253 -631
rect -219 -665 -213 -631
rect -259 -703 -213 -665
rect -259 -737 -253 -703
rect -219 -737 -213 -703
rect -259 -775 -213 -737
rect -259 -809 -253 -775
rect -219 -809 -213 -775
rect -259 -847 -213 -809
rect -259 -881 -253 -847
rect -219 -881 -213 -847
rect -259 -919 -213 -881
rect -259 -953 -253 -919
rect -219 -953 -213 -919
rect -259 -991 -213 -953
rect -259 -1025 -253 -991
rect -219 -1025 -213 -991
rect -259 -1063 -213 -1025
rect -259 -1097 -253 -1063
rect -219 -1097 -213 -1063
rect -259 -1135 -213 -1097
rect -259 -1169 -253 -1135
rect -219 -1169 -213 -1135
rect -259 -1207 -213 -1169
rect -259 -1241 -253 -1207
rect -219 -1241 -213 -1207
rect -259 -1279 -213 -1241
rect -259 -1313 -253 -1279
rect -219 -1313 -213 -1279
rect -259 -1351 -213 -1313
rect -259 -1385 -253 -1351
rect -219 -1385 -213 -1351
rect -259 -1423 -213 -1385
rect -259 -1457 -253 -1423
rect -219 -1457 -213 -1423
rect -259 -1500 -213 -1457
rect -141 1457 -95 1500
rect -141 1423 -135 1457
rect -101 1423 -95 1457
rect -141 1385 -95 1423
rect -141 1351 -135 1385
rect -101 1351 -95 1385
rect -141 1313 -95 1351
rect -141 1279 -135 1313
rect -101 1279 -95 1313
rect -141 1241 -95 1279
rect -141 1207 -135 1241
rect -101 1207 -95 1241
rect -141 1169 -95 1207
rect -141 1135 -135 1169
rect -101 1135 -95 1169
rect -141 1097 -95 1135
rect -141 1063 -135 1097
rect -101 1063 -95 1097
rect -141 1025 -95 1063
rect -141 991 -135 1025
rect -101 991 -95 1025
rect -141 953 -95 991
rect -141 919 -135 953
rect -101 919 -95 953
rect -141 881 -95 919
rect -141 847 -135 881
rect -101 847 -95 881
rect -141 809 -95 847
rect -141 775 -135 809
rect -101 775 -95 809
rect -141 737 -95 775
rect -141 703 -135 737
rect -101 703 -95 737
rect -141 665 -95 703
rect -141 631 -135 665
rect -101 631 -95 665
rect -141 593 -95 631
rect -141 559 -135 593
rect -101 559 -95 593
rect -141 521 -95 559
rect -141 487 -135 521
rect -101 487 -95 521
rect -141 449 -95 487
rect -141 415 -135 449
rect -101 415 -95 449
rect -141 377 -95 415
rect -141 343 -135 377
rect -101 343 -95 377
rect -141 305 -95 343
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -343 -95 -305
rect -141 -377 -135 -343
rect -101 -377 -95 -343
rect -141 -415 -95 -377
rect -141 -449 -135 -415
rect -101 -449 -95 -415
rect -141 -487 -95 -449
rect -141 -521 -135 -487
rect -101 -521 -95 -487
rect -141 -559 -95 -521
rect -141 -593 -135 -559
rect -101 -593 -95 -559
rect -141 -631 -95 -593
rect -141 -665 -135 -631
rect -101 -665 -95 -631
rect -141 -703 -95 -665
rect -141 -737 -135 -703
rect -101 -737 -95 -703
rect -141 -775 -95 -737
rect -141 -809 -135 -775
rect -101 -809 -95 -775
rect -141 -847 -95 -809
rect -141 -881 -135 -847
rect -101 -881 -95 -847
rect -141 -919 -95 -881
rect -141 -953 -135 -919
rect -101 -953 -95 -919
rect -141 -991 -95 -953
rect -141 -1025 -135 -991
rect -101 -1025 -95 -991
rect -141 -1063 -95 -1025
rect -141 -1097 -135 -1063
rect -101 -1097 -95 -1063
rect -141 -1135 -95 -1097
rect -141 -1169 -135 -1135
rect -101 -1169 -95 -1135
rect -141 -1207 -95 -1169
rect -141 -1241 -135 -1207
rect -101 -1241 -95 -1207
rect -141 -1279 -95 -1241
rect -141 -1313 -135 -1279
rect -101 -1313 -95 -1279
rect -141 -1351 -95 -1313
rect -141 -1385 -135 -1351
rect -101 -1385 -95 -1351
rect -141 -1423 -95 -1385
rect -141 -1457 -135 -1423
rect -101 -1457 -95 -1423
rect -141 -1500 -95 -1457
rect -23 1457 23 1500
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1500 23 -1457
rect 95 1457 141 1500
rect 95 1423 101 1457
rect 135 1423 141 1457
rect 95 1385 141 1423
rect 95 1351 101 1385
rect 135 1351 141 1385
rect 95 1313 141 1351
rect 95 1279 101 1313
rect 135 1279 141 1313
rect 95 1241 141 1279
rect 95 1207 101 1241
rect 135 1207 141 1241
rect 95 1169 141 1207
rect 95 1135 101 1169
rect 135 1135 141 1169
rect 95 1097 141 1135
rect 95 1063 101 1097
rect 135 1063 141 1097
rect 95 1025 141 1063
rect 95 991 101 1025
rect 135 991 141 1025
rect 95 953 141 991
rect 95 919 101 953
rect 135 919 141 953
rect 95 881 141 919
rect 95 847 101 881
rect 135 847 141 881
rect 95 809 141 847
rect 95 775 101 809
rect 135 775 141 809
rect 95 737 141 775
rect 95 703 101 737
rect 135 703 141 737
rect 95 665 141 703
rect 95 631 101 665
rect 135 631 141 665
rect 95 593 141 631
rect 95 559 101 593
rect 135 559 141 593
rect 95 521 141 559
rect 95 487 101 521
rect 135 487 141 521
rect 95 449 141 487
rect 95 415 101 449
rect 135 415 141 449
rect 95 377 141 415
rect 95 343 101 377
rect 135 343 141 377
rect 95 305 141 343
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -343 141 -305
rect 95 -377 101 -343
rect 135 -377 141 -343
rect 95 -415 141 -377
rect 95 -449 101 -415
rect 135 -449 141 -415
rect 95 -487 141 -449
rect 95 -521 101 -487
rect 135 -521 141 -487
rect 95 -559 141 -521
rect 95 -593 101 -559
rect 135 -593 141 -559
rect 95 -631 141 -593
rect 95 -665 101 -631
rect 135 -665 141 -631
rect 95 -703 141 -665
rect 95 -737 101 -703
rect 135 -737 141 -703
rect 95 -775 141 -737
rect 95 -809 101 -775
rect 135 -809 141 -775
rect 95 -847 141 -809
rect 95 -881 101 -847
rect 135 -881 141 -847
rect 95 -919 141 -881
rect 95 -953 101 -919
rect 135 -953 141 -919
rect 95 -991 141 -953
rect 95 -1025 101 -991
rect 135 -1025 141 -991
rect 95 -1063 141 -1025
rect 95 -1097 101 -1063
rect 135 -1097 141 -1063
rect 95 -1135 141 -1097
rect 95 -1169 101 -1135
rect 135 -1169 141 -1135
rect 95 -1207 141 -1169
rect 95 -1241 101 -1207
rect 135 -1241 141 -1207
rect 95 -1279 141 -1241
rect 95 -1313 101 -1279
rect 135 -1313 141 -1279
rect 95 -1351 141 -1313
rect 95 -1385 101 -1351
rect 135 -1385 141 -1351
rect 95 -1423 141 -1385
rect 95 -1457 101 -1423
rect 135 -1457 141 -1423
rect 95 -1500 141 -1457
rect 213 1457 259 1500
rect 213 1423 219 1457
rect 253 1423 259 1457
rect 213 1385 259 1423
rect 213 1351 219 1385
rect 253 1351 259 1385
rect 213 1313 259 1351
rect 213 1279 219 1313
rect 253 1279 259 1313
rect 213 1241 259 1279
rect 213 1207 219 1241
rect 253 1207 259 1241
rect 213 1169 259 1207
rect 213 1135 219 1169
rect 253 1135 259 1169
rect 213 1097 259 1135
rect 213 1063 219 1097
rect 253 1063 259 1097
rect 213 1025 259 1063
rect 213 991 219 1025
rect 253 991 259 1025
rect 213 953 259 991
rect 213 919 219 953
rect 253 919 259 953
rect 213 881 259 919
rect 213 847 219 881
rect 253 847 259 881
rect 213 809 259 847
rect 213 775 219 809
rect 253 775 259 809
rect 213 737 259 775
rect 213 703 219 737
rect 253 703 259 737
rect 213 665 259 703
rect 213 631 219 665
rect 253 631 259 665
rect 213 593 259 631
rect 213 559 219 593
rect 253 559 259 593
rect 213 521 259 559
rect 213 487 219 521
rect 253 487 259 521
rect 213 449 259 487
rect 213 415 219 449
rect 253 415 259 449
rect 213 377 259 415
rect 213 343 219 377
rect 253 343 259 377
rect 213 305 259 343
rect 213 271 219 305
rect 253 271 259 305
rect 213 233 259 271
rect 213 199 219 233
rect 253 199 259 233
rect 213 161 259 199
rect 213 127 219 161
rect 253 127 259 161
rect 213 89 259 127
rect 213 55 219 89
rect 253 55 259 89
rect 213 17 259 55
rect 213 -17 219 17
rect 253 -17 259 17
rect 213 -55 259 -17
rect 213 -89 219 -55
rect 253 -89 259 -55
rect 213 -127 259 -89
rect 213 -161 219 -127
rect 253 -161 259 -127
rect 213 -199 259 -161
rect 213 -233 219 -199
rect 253 -233 259 -199
rect 213 -271 259 -233
rect 213 -305 219 -271
rect 253 -305 259 -271
rect 213 -343 259 -305
rect 213 -377 219 -343
rect 253 -377 259 -343
rect 213 -415 259 -377
rect 213 -449 219 -415
rect 253 -449 259 -415
rect 213 -487 259 -449
rect 213 -521 219 -487
rect 253 -521 259 -487
rect 213 -559 259 -521
rect 213 -593 219 -559
rect 253 -593 259 -559
rect 213 -631 259 -593
rect 213 -665 219 -631
rect 253 -665 259 -631
rect 213 -703 259 -665
rect 213 -737 219 -703
rect 253 -737 259 -703
rect 213 -775 259 -737
rect 213 -809 219 -775
rect 253 -809 259 -775
rect 213 -847 259 -809
rect 213 -881 219 -847
rect 253 -881 259 -847
rect 213 -919 259 -881
rect 213 -953 219 -919
rect 253 -953 259 -919
rect 213 -991 259 -953
rect 213 -1025 219 -991
rect 253 -1025 259 -991
rect 213 -1063 259 -1025
rect 213 -1097 219 -1063
rect 253 -1097 259 -1063
rect 213 -1135 259 -1097
rect 213 -1169 219 -1135
rect 253 -1169 259 -1135
rect 213 -1207 259 -1169
rect 213 -1241 219 -1207
rect 253 -1241 259 -1207
rect 213 -1279 259 -1241
rect 213 -1313 219 -1279
rect 253 -1313 259 -1279
rect 213 -1351 259 -1313
rect 213 -1385 219 -1351
rect 253 -1385 259 -1351
rect 213 -1423 259 -1385
rect 213 -1457 219 -1423
rect 253 -1457 259 -1423
rect 213 -1500 259 -1457
rect -206 -1547 -148 -1541
rect -206 -1581 -194 -1547
rect -160 -1581 -148 -1547
rect -206 -1587 -148 -1581
rect -88 -1547 -30 -1541
rect -88 -1581 -76 -1547
rect -42 -1581 -30 -1547
rect -88 -1587 -30 -1581
rect 30 -1547 88 -1541
rect 30 -1581 42 -1547
rect 76 -1581 88 -1547
rect 30 -1587 88 -1581
rect 148 -1547 206 -1541
rect 148 -1581 160 -1547
rect 194 -1581 206 -1547
rect 148 -1587 206 -1581
<< properties >>
string FIXED_BBOX -350 -1666 350 1666
<< end >>
