//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: maskmul
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Jan 15 17:23:49 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

module maskmul_top_formal_verification (
input [0:0] am_0_,
input [0:0] am_1_,
input [0:0] bm_0_,
input [0:0] bm_1_,
input [0:0] ma_0_,
input [0:0] ma_1_,
input [0:0] mb_0_,
input [0:0] mb_1_,
input [0:0] mq_0_,
input [0:0] mq_1_,
input [0:0] reset,
input [0:0] clk,
output [0:0] qm_0_,
output [0:0] qm_1_);

// ----- Local wires for FPGA fabric -----
wire [0:63] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] prog_clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;
wire [0:0] clk_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		.prog_clk(prog_clk_fm[0]),
		.set(set_fm[0]),
		.reset(reset_fm[0]),
		.clk(clk_fm[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD_fm[0:63]),
		.ccff_head(ccff_head_fm[0]),
		.ccff_tail(ccff_tail_fm[0]));

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = reset[0];
	assign clk_fm[0] = clk[0];
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input am_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[35] -----
	assign gfpga_pad_GPIO_PAD_fm[35] = am_0_[0];

// ----- Blif Benchmark input am_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[41] -----
	assign gfpga_pad_GPIO_PAD_fm[41] = am_1_[0];

// ----- Blif Benchmark input bm_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[34] -----
	assign gfpga_pad_GPIO_PAD_fm[34] = bm_0_[0];

// ----- Blif Benchmark input bm_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[42] -----
	assign gfpga_pad_GPIO_PAD_fm[42] = bm_1_[0];

// ----- Blif Benchmark input ma_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[28] -----
	assign gfpga_pad_GPIO_PAD_fm[28] = ma_0_[0];

// ----- Blif Benchmark input ma_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[55] -----
	assign gfpga_pad_GPIO_PAD_fm[55] = ma_1_[0];

// ----- Blif Benchmark input mb_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[33] -----
	assign gfpga_pad_GPIO_PAD_fm[33] = mb_0_[0];

// ----- Blif Benchmark input mb_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[40] -----
	assign gfpga_pad_GPIO_PAD_fm[40] = mb_1_[0];

// ----- Blif Benchmark input mq_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[47] -----
	assign gfpga_pad_GPIO_PAD_fm[47] = mq_0_[0];

// ----- Blif Benchmark input mq_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[31] -----
	assign gfpga_pad_GPIO_PAD_fm[31] = mq_1_[0];

// ----- Blif Benchmark input reset is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[44] -----
	assign gfpga_pad_GPIO_PAD_fm[44] = reset[0];

// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[53] -----
	assign gfpga_pad_GPIO_PAD_fm[53] = clk[0];

// ----- Blif Benchmark output qm_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[48] -----
	assign qm_0_[0] = gfpga_pad_GPIO_PAD_fm[48];

// ----- Blif Benchmark output qm_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[26] -----
	assign qm_1_[0] = gfpga_pad_GPIO_PAD_fm[26];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[32] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[50] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[54] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[56] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[62] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[63] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin deposit bitstream to configuration memories -----
initial begin
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0001001001001000);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1110110110110111);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0110011001100110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1001100110011001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0001001001001000);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1110110110110111);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0000000010010110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1111111101101001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3], 4'b0010);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3], 4'b1101);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3], 4'b1101);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3], 4'b0010);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3], 4'b1001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3], 4'b0110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3], 4'b0011);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3], 4'b1100);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3], 4'b1011);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3], 4'b0100);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3], 4'b0011);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3], 4'b1100);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3], 4'b1011);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3], 4'b0100);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3], 4'b1101);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3], 4'b0010);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3], 4'b1100);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3], 4'b0011);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3], 4'b0111);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3], 4'b1000);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3], 4'b0001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3], 4'b1110);
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0110011001100110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1001100110011001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0001001001001000);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1110110110110111);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b1001101001101010);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b0110010110010101);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], 16'b0001001000010010);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], 16'b1110110111101101);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3], 4'b1011);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3], 4'b0100);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3], 4'b0001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3], 4'b1110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3], 4'b1011);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3], 4'b0100);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3], 4'b1110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3], 4'b0001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3], 4'b0001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3], 4'b1110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3], 4'b0011);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3], 4'b1100);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3], 4'b1110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3], 4'b0001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3], 4'b1001);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3], 4'b0110);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3], 4'b0111);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3], 4'b1000);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3], 4'b1100);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3], 4'b0011);
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:3], 4'b0001);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:3], 4'b1110);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:3], 4'b0101);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:3], 4'b1010);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:3], 4'b0010);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:3], 4'b1101);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3], 4'b0101);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:3], 4'b1010);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3], 4'b0001);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:3], 4'b1110);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3], 4'b0010);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3], 4'b1101);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3], 4'b0010);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:3], 4'b1101);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3], 4'b0100);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:3], 4'b1011);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:3], 4'b0011);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:3], 4'b1100);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3], 4'b0110);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:3], 4'b1001);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_3.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_7.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_7.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:2], 3'b011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:2], 3'b100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:2], 3'b110);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:2], 3'b001);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:2], 3'b101);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:2], 3'b010);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:2], 3'b101);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:2], 3'b011);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:2], 3'b100);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_out[0:2], 3'b101);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_outb[0:2], 3'b010);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b1}});
end
// ----- End deposit bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for maskmul_top_formal_verification -----

