magic
tech sky130A
magscale 1 2
timestamp 1752660100
<< pwell >>
rect -201 -742 201 742
<< psubdiff >>
rect -165 672 -69 706
rect 69 672 165 706
rect -165 610 -131 672
rect 131 610 165 672
rect -165 -672 -131 -610
rect 131 -672 165 -610
rect -165 -706 -69 -672
rect 69 -706 165 -672
<< psubdiffcont >>
rect -69 672 69 706
rect -165 -610 -131 610
rect 131 -610 165 610
rect -69 -706 69 -672
<< xpolycontact >>
rect -35 144 35 576
rect -35 -576 35 -144
<< xpolyres >>
rect -35 -144 35 144
<< locali >>
rect -165 672 -69 706
rect 69 672 165 706
rect -165 610 -131 672
rect 131 610 165 672
rect -165 -672 -131 -610
rect 131 -672 165 -610
rect -165 -706 -69 -672
rect 69 -706 165 -672
<< viali >>
rect -19 161 19 558
rect -19 -558 19 -161
<< metal1 >>
rect -25 558 25 570
rect -25 161 -19 558
rect 19 161 25 558
rect -25 149 25 161
rect -25 -161 25 -149
rect -25 -558 -19 -161
rect 19 -558 25 -161
rect -25 -570 25 -558
<< properties >>
string FIXED_BBOX -148 -689 148 689
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.6 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 10.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
