magic
tech sky130A
magscale 1 2
timestamp 1757256347
<< pwell >>
rect -280 -327 280 327
<< mvnmos >>
rect -50 -131 50 69
<< mvndiff >>
rect -108 57 -50 69
rect -108 -119 -96 57
rect -62 -119 -50 57
rect -108 -131 -50 -119
rect 50 57 108 69
rect 50 -119 62 57
rect 96 -119 108 57
rect 50 -131 108 -119
<< mvndiffc >>
rect -96 -119 -62 57
rect 62 -119 96 57
<< mvpsubdiff >>
rect -244 279 244 291
rect -244 245 -136 279
rect 136 245 244 279
rect -244 233 244 245
rect -244 183 -186 233
rect -244 -183 -232 183
rect -198 -183 -186 183
rect 186 183 244 233
rect -244 -233 -186 -183
rect 186 -183 198 183
rect 232 -183 244 183
rect 186 -233 244 -183
rect -244 -245 244 -233
rect -244 -279 -136 -245
rect 136 -279 244 -245
rect -244 -291 244 -279
<< mvpsubdiffcont >>
rect -136 245 136 279
rect -232 -183 -198 183
rect 198 -183 232 183
rect -136 -279 136 -245
<< poly >>
rect -50 141 50 157
rect -50 107 -34 141
rect 34 107 50 141
rect -50 69 50 107
rect -50 -157 50 -131
<< polycont >>
rect -34 107 34 141
<< locali >>
rect -232 245 -136 279
rect 136 245 232 279
rect -232 183 -198 245
rect 198 183 232 245
rect -50 107 -34 141
rect 34 107 50 141
rect -96 57 -62 73
rect -96 -135 -62 -119
rect 62 57 96 73
rect 62 -135 96 -119
rect -232 -245 -198 -183
rect 198 -245 232 -183
rect -232 -279 -136 -245
rect 136 -279 232 -245
<< viali >>
rect -34 107 34 141
rect -96 -119 -62 57
rect 62 -119 96 57
<< metal1 >>
rect -46 141 46 147
rect -46 107 -34 141
rect 34 107 46 141
rect -46 101 46 107
rect -102 57 -56 69
rect -102 -119 -96 57
rect -62 -119 -56 57
rect -102 -131 -56 -119
rect 56 57 102 69
rect 56 -119 62 57
rect 96 -119 102 57
rect 56 -131 102 -119
<< labels >>
rlabel mvpsubdiffcont 0 -262 0 -262 0 B
port 1 nsew
rlabel mvndiffc -79 -31 -79 -31 0 D
port 2 nsew
rlabel mvndiffc 79 -31 79 -31 0 S
port 3 nsew
rlabel polycont 0 124 0 124 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -215 -262 215 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
