magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -365 881 -307 887
rect -173 881 -115 887
rect 19 881 77 887
rect 211 881 269 887
rect 403 881 461 887
rect -365 847 -353 881
rect -173 847 -161 881
rect 19 847 31 881
rect 211 847 223 881
rect 403 847 415 881
rect -365 841 -307 847
rect -173 841 -115 847
rect 19 841 77 847
rect 211 841 269 847
rect 403 841 461 847
rect -461 -847 -403 -841
rect -269 -847 -211 -841
rect -77 -847 -19 -841
rect 115 -847 173 -841
rect 307 -847 365 -841
rect -461 -881 -449 -847
rect -269 -881 -257 -847
rect -77 -881 -65 -847
rect 115 -881 127 -847
rect 307 -881 319 -847
rect -461 -887 -403 -881
rect -269 -887 -211 -881
rect -77 -887 -19 -881
rect 115 -887 173 -881
rect 307 -887 365 -881
<< nwell >>
rect -647 -1019 647 1019
<< pmos >>
rect -447 -800 -417 800
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
rect 417 -800 447 800
<< pdiff >>
rect -509 765 -447 800
rect -509 731 -497 765
rect -463 731 -447 765
rect -509 697 -447 731
rect -509 663 -497 697
rect -463 663 -447 697
rect -509 629 -447 663
rect -509 595 -497 629
rect -463 595 -447 629
rect -509 561 -447 595
rect -509 527 -497 561
rect -463 527 -447 561
rect -509 493 -447 527
rect -509 459 -497 493
rect -463 459 -447 493
rect -509 425 -447 459
rect -509 391 -497 425
rect -463 391 -447 425
rect -509 357 -447 391
rect -509 323 -497 357
rect -463 323 -447 357
rect -509 289 -447 323
rect -509 255 -497 289
rect -463 255 -447 289
rect -509 221 -447 255
rect -509 187 -497 221
rect -463 187 -447 221
rect -509 153 -447 187
rect -509 119 -497 153
rect -463 119 -447 153
rect -509 85 -447 119
rect -509 51 -497 85
rect -463 51 -447 85
rect -509 17 -447 51
rect -509 -17 -497 17
rect -463 -17 -447 17
rect -509 -51 -447 -17
rect -509 -85 -497 -51
rect -463 -85 -447 -51
rect -509 -119 -447 -85
rect -509 -153 -497 -119
rect -463 -153 -447 -119
rect -509 -187 -447 -153
rect -509 -221 -497 -187
rect -463 -221 -447 -187
rect -509 -255 -447 -221
rect -509 -289 -497 -255
rect -463 -289 -447 -255
rect -509 -323 -447 -289
rect -509 -357 -497 -323
rect -463 -357 -447 -323
rect -509 -391 -447 -357
rect -509 -425 -497 -391
rect -463 -425 -447 -391
rect -509 -459 -447 -425
rect -509 -493 -497 -459
rect -463 -493 -447 -459
rect -509 -527 -447 -493
rect -509 -561 -497 -527
rect -463 -561 -447 -527
rect -509 -595 -447 -561
rect -509 -629 -497 -595
rect -463 -629 -447 -595
rect -509 -663 -447 -629
rect -509 -697 -497 -663
rect -463 -697 -447 -663
rect -509 -731 -447 -697
rect -509 -765 -497 -731
rect -463 -765 -447 -731
rect -509 -800 -447 -765
rect -417 765 -351 800
rect -417 731 -401 765
rect -367 731 -351 765
rect -417 697 -351 731
rect -417 663 -401 697
rect -367 663 -351 697
rect -417 629 -351 663
rect -417 595 -401 629
rect -367 595 -351 629
rect -417 561 -351 595
rect -417 527 -401 561
rect -367 527 -351 561
rect -417 493 -351 527
rect -417 459 -401 493
rect -367 459 -351 493
rect -417 425 -351 459
rect -417 391 -401 425
rect -367 391 -351 425
rect -417 357 -351 391
rect -417 323 -401 357
rect -367 323 -351 357
rect -417 289 -351 323
rect -417 255 -401 289
rect -367 255 -351 289
rect -417 221 -351 255
rect -417 187 -401 221
rect -367 187 -351 221
rect -417 153 -351 187
rect -417 119 -401 153
rect -367 119 -351 153
rect -417 85 -351 119
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -119 -351 -85
rect -417 -153 -401 -119
rect -367 -153 -351 -119
rect -417 -187 -351 -153
rect -417 -221 -401 -187
rect -367 -221 -351 -187
rect -417 -255 -351 -221
rect -417 -289 -401 -255
rect -367 -289 -351 -255
rect -417 -323 -351 -289
rect -417 -357 -401 -323
rect -367 -357 -351 -323
rect -417 -391 -351 -357
rect -417 -425 -401 -391
rect -367 -425 -351 -391
rect -417 -459 -351 -425
rect -417 -493 -401 -459
rect -367 -493 -351 -459
rect -417 -527 -351 -493
rect -417 -561 -401 -527
rect -367 -561 -351 -527
rect -417 -595 -351 -561
rect -417 -629 -401 -595
rect -367 -629 -351 -595
rect -417 -663 -351 -629
rect -417 -697 -401 -663
rect -367 -697 -351 -663
rect -417 -731 -351 -697
rect -417 -765 -401 -731
rect -367 -765 -351 -731
rect -417 -800 -351 -765
rect -321 765 -255 800
rect -321 731 -305 765
rect -271 731 -255 765
rect -321 697 -255 731
rect -321 663 -305 697
rect -271 663 -255 697
rect -321 629 -255 663
rect -321 595 -305 629
rect -271 595 -255 629
rect -321 561 -255 595
rect -321 527 -305 561
rect -271 527 -255 561
rect -321 493 -255 527
rect -321 459 -305 493
rect -271 459 -255 493
rect -321 425 -255 459
rect -321 391 -305 425
rect -271 391 -255 425
rect -321 357 -255 391
rect -321 323 -305 357
rect -271 323 -255 357
rect -321 289 -255 323
rect -321 255 -305 289
rect -271 255 -255 289
rect -321 221 -255 255
rect -321 187 -305 221
rect -271 187 -255 221
rect -321 153 -255 187
rect -321 119 -305 153
rect -271 119 -255 153
rect -321 85 -255 119
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -119 -255 -85
rect -321 -153 -305 -119
rect -271 -153 -255 -119
rect -321 -187 -255 -153
rect -321 -221 -305 -187
rect -271 -221 -255 -187
rect -321 -255 -255 -221
rect -321 -289 -305 -255
rect -271 -289 -255 -255
rect -321 -323 -255 -289
rect -321 -357 -305 -323
rect -271 -357 -255 -323
rect -321 -391 -255 -357
rect -321 -425 -305 -391
rect -271 -425 -255 -391
rect -321 -459 -255 -425
rect -321 -493 -305 -459
rect -271 -493 -255 -459
rect -321 -527 -255 -493
rect -321 -561 -305 -527
rect -271 -561 -255 -527
rect -321 -595 -255 -561
rect -321 -629 -305 -595
rect -271 -629 -255 -595
rect -321 -663 -255 -629
rect -321 -697 -305 -663
rect -271 -697 -255 -663
rect -321 -731 -255 -697
rect -321 -765 -305 -731
rect -271 -765 -255 -731
rect -321 -800 -255 -765
rect -225 765 -159 800
rect -225 731 -209 765
rect -175 731 -159 765
rect -225 697 -159 731
rect -225 663 -209 697
rect -175 663 -159 697
rect -225 629 -159 663
rect -225 595 -209 629
rect -175 595 -159 629
rect -225 561 -159 595
rect -225 527 -209 561
rect -175 527 -159 561
rect -225 493 -159 527
rect -225 459 -209 493
rect -175 459 -159 493
rect -225 425 -159 459
rect -225 391 -209 425
rect -175 391 -159 425
rect -225 357 -159 391
rect -225 323 -209 357
rect -175 323 -159 357
rect -225 289 -159 323
rect -225 255 -209 289
rect -175 255 -159 289
rect -225 221 -159 255
rect -225 187 -209 221
rect -175 187 -159 221
rect -225 153 -159 187
rect -225 119 -209 153
rect -175 119 -159 153
rect -225 85 -159 119
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -119 -159 -85
rect -225 -153 -209 -119
rect -175 -153 -159 -119
rect -225 -187 -159 -153
rect -225 -221 -209 -187
rect -175 -221 -159 -187
rect -225 -255 -159 -221
rect -225 -289 -209 -255
rect -175 -289 -159 -255
rect -225 -323 -159 -289
rect -225 -357 -209 -323
rect -175 -357 -159 -323
rect -225 -391 -159 -357
rect -225 -425 -209 -391
rect -175 -425 -159 -391
rect -225 -459 -159 -425
rect -225 -493 -209 -459
rect -175 -493 -159 -459
rect -225 -527 -159 -493
rect -225 -561 -209 -527
rect -175 -561 -159 -527
rect -225 -595 -159 -561
rect -225 -629 -209 -595
rect -175 -629 -159 -595
rect -225 -663 -159 -629
rect -225 -697 -209 -663
rect -175 -697 -159 -663
rect -225 -731 -159 -697
rect -225 -765 -209 -731
rect -175 -765 -159 -731
rect -225 -800 -159 -765
rect -129 765 -63 800
rect -129 731 -113 765
rect -79 731 -63 765
rect -129 697 -63 731
rect -129 663 -113 697
rect -79 663 -63 697
rect -129 629 -63 663
rect -129 595 -113 629
rect -79 595 -63 629
rect -129 561 -63 595
rect -129 527 -113 561
rect -79 527 -63 561
rect -129 493 -63 527
rect -129 459 -113 493
rect -79 459 -63 493
rect -129 425 -63 459
rect -129 391 -113 425
rect -79 391 -63 425
rect -129 357 -63 391
rect -129 323 -113 357
rect -79 323 -63 357
rect -129 289 -63 323
rect -129 255 -113 289
rect -79 255 -63 289
rect -129 221 -63 255
rect -129 187 -113 221
rect -79 187 -63 221
rect -129 153 -63 187
rect -129 119 -113 153
rect -79 119 -63 153
rect -129 85 -63 119
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -119 -63 -85
rect -129 -153 -113 -119
rect -79 -153 -63 -119
rect -129 -187 -63 -153
rect -129 -221 -113 -187
rect -79 -221 -63 -187
rect -129 -255 -63 -221
rect -129 -289 -113 -255
rect -79 -289 -63 -255
rect -129 -323 -63 -289
rect -129 -357 -113 -323
rect -79 -357 -63 -323
rect -129 -391 -63 -357
rect -129 -425 -113 -391
rect -79 -425 -63 -391
rect -129 -459 -63 -425
rect -129 -493 -113 -459
rect -79 -493 -63 -459
rect -129 -527 -63 -493
rect -129 -561 -113 -527
rect -79 -561 -63 -527
rect -129 -595 -63 -561
rect -129 -629 -113 -595
rect -79 -629 -63 -595
rect -129 -663 -63 -629
rect -129 -697 -113 -663
rect -79 -697 -63 -663
rect -129 -731 -63 -697
rect -129 -765 -113 -731
rect -79 -765 -63 -731
rect -129 -800 -63 -765
rect -33 765 33 800
rect -33 731 -17 765
rect 17 731 33 765
rect -33 697 33 731
rect -33 663 -17 697
rect 17 663 33 697
rect -33 629 33 663
rect -33 595 -17 629
rect 17 595 33 629
rect -33 561 33 595
rect -33 527 -17 561
rect 17 527 33 561
rect -33 493 33 527
rect -33 459 -17 493
rect 17 459 33 493
rect -33 425 33 459
rect -33 391 -17 425
rect 17 391 33 425
rect -33 357 33 391
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -391 33 -357
rect -33 -425 -17 -391
rect 17 -425 33 -391
rect -33 -459 33 -425
rect -33 -493 -17 -459
rect 17 -493 33 -459
rect -33 -527 33 -493
rect -33 -561 -17 -527
rect 17 -561 33 -527
rect -33 -595 33 -561
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -663 33 -629
rect -33 -697 -17 -663
rect 17 -697 33 -663
rect -33 -731 33 -697
rect -33 -765 -17 -731
rect 17 -765 33 -731
rect -33 -800 33 -765
rect 63 765 129 800
rect 63 731 79 765
rect 113 731 129 765
rect 63 697 129 731
rect 63 663 79 697
rect 113 663 129 697
rect 63 629 129 663
rect 63 595 79 629
rect 113 595 129 629
rect 63 561 129 595
rect 63 527 79 561
rect 113 527 129 561
rect 63 493 129 527
rect 63 459 79 493
rect 113 459 129 493
rect 63 425 129 459
rect 63 391 79 425
rect 113 391 129 425
rect 63 357 129 391
rect 63 323 79 357
rect 113 323 129 357
rect 63 289 129 323
rect 63 255 79 289
rect 113 255 129 289
rect 63 221 129 255
rect 63 187 79 221
rect 113 187 129 221
rect 63 153 129 187
rect 63 119 79 153
rect 113 119 129 153
rect 63 85 129 119
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -119 129 -85
rect 63 -153 79 -119
rect 113 -153 129 -119
rect 63 -187 129 -153
rect 63 -221 79 -187
rect 113 -221 129 -187
rect 63 -255 129 -221
rect 63 -289 79 -255
rect 113 -289 129 -255
rect 63 -323 129 -289
rect 63 -357 79 -323
rect 113 -357 129 -323
rect 63 -391 129 -357
rect 63 -425 79 -391
rect 113 -425 129 -391
rect 63 -459 129 -425
rect 63 -493 79 -459
rect 113 -493 129 -459
rect 63 -527 129 -493
rect 63 -561 79 -527
rect 113 -561 129 -527
rect 63 -595 129 -561
rect 63 -629 79 -595
rect 113 -629 129 -595
rect 63 -663 129 -629
rect 63 -697 79 -663
rect 113 -697 129 -663
rect 63 -731 129 -697
rect 63 -765 79 -731
rect 113 -765 129 -731
rect 63 -800 129 -765
rect 159 765 225 800
rect 159 731 175 765
rect 209 731 225 765
rect 159 697 225 731
rect 159 663 175 697
rect 209 663 225 697
rect 159 629 225 663
rect 159 595 175 629
rect 209 595 225 629
rect 159 561 225 595
rect 159 527 175 561
rect 209 527 225 561
rect 159 493 225 527
rect 159 459 175 493
rect 209 459 225 493
rect 159 425 225 459
rect 159 391 175 425
rect 209 391 225 425
rect 159 357 225 391
rect 159 323 175 357
rect 209 323 225 357
rect 159 289 225 323
rect 159 255 175 289
rect 209 255 225 289
rect 159 221 225 255
rect 159 187 175 221
rect 209 187 225 221
rect 159 153 225 187
rect 159 119 175 153
rect 209 119 225 153
rect 159 85 225 119
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -119 225 -85
rect 159 -153 175 -119
rect 209 -153 225 -119
rect 159 -187 225 -153
rect 159 -221 175 -187
rect 209 -221 225 -187
rect 159 -255 225 -221
rect 159 -289 175 -255
rect 209 -289 225 -255
rect 159 -323 225 -289
rect 159 -357 175 -323
rect 209 -357 225 -323
rect 159 -391 225 -357
rect 159 -425 175 -391
rect 209 -425 225 -391
rect 159 -459 225 -425
rect 159 -493 175 -459
rect 209 -493 225 -459
rect 159 -527 225 -493
rect 159 -561 175 -527
rect 209 -561 225 -527
rect 159 -595 225 -561
rect 159 -629 175 -595
rect 209 -629 225 -595
rect 159 -663 225 -629
rect 159 -697 175 -663
rect 209 -697 225 -663
rect 159 -731 225 -697
rect 159 -765 175 -731
rect 209 -765 225 -731
rect 159 -800 225 -765
rect 255 765 321 800
rect 255 731 271 765
rect 305 731 321 765
rect 255 697 321 731
rect 255 663 271 697
rect 305 663 321 697
rect 255 629 321 663
rect 255 595 271 629
rect 305 595 321 629
rect 255 561 321 595
rect 255 527 271 561
rect 305 527 321 561
rect 255 493 321 527
rect 255 459 271 493
rect 305 459 321 493
rect 255 425 321 459
rect 255 391 271 425
rect 305 391 321 425
rect 255 357 321 391
rect 255 323 271 357
rect 305 323 321 357
rect 255 289 321 323
rect 255 255 271 289
rect 305 255 321 289
rect 255 221 321 255
rect 255 187 271 221
rect 305 187 321 221
rect 255 153 321 187
rect 255 119 271 153
rect 305 119 321 153
rect 255 85 321 119
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -119 321 -85
rect 255 -153 271 -119
rect 305 -153 321 -119
rect 255 -187 321 -153
rect 255 -221 271 -187
rect 305 -221 321 -187
rect 255 -255 321 -221
rect 255 -289 271 -255
rect 305 -289 321 -255
rect 255 -323 321 -289
rect 255 -357 271 -323
rect 305 -357 321 -323
rect 255 -391 321 -357
rect 255 -425 271 -391
rect 305 -425 321 -391
rect 255 -459 321 -425
rect 255 -493 271 -459
rect 305 -493 321 -459
rect 255 -527 321 -493
rect 255 -561 271 -527
rect 305 -561 321 -527
rect 255 -595 321 -561
rect 255 -629 271 -595
rect 305 -629 321 -595
rect 255 -663 321 -629
rect 255 -697 271 -663
rect 305 -697 321 -663
rect 255 -731 321 -697
rect 255 -765 271 -731
rect 305 -765 321 -731
rect 255 -800 321 -765
rect 351 765 417 800
rect 351 731 367 765
rect 401 731 417 765
rect 351 697 417 731
rect 351 663 367 697
rect 401 663 417 697
rect 351 629 417 663
rect 351 595 367 629
rect 401 595 417 629
rect 351 561 417 595
rect 351 527 367 561
rect 401 527 417 561
rect 351 493 417 527
rect 351 459 367 493
rect 401 459 417 493
rect 351 425 417 459
rect 351 391 367 425
rect 401 391 417 425
rect 351 357 417 391
rect 351 323 367 357
rect 401 323 417 357
rect 351 289 417 323
rect 351 255 367 289
rect 401 255 417 289
rect 351 221 417 255
rect 351 187 367 221
rect 401 187 417 221
rect 351 153 417 187
rect 351 119 367 153
rect 401 119 417 153
rect 351 85 417 119
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -119 417 -85
rect 351 -153 367 -119
rect 401 -153 417 -119
rect 351 -187 417 -153
rect 351 -221 367 -187
rect 401 -221 417 -187
rect 351 -255 417 -221
rect 351 -289 367 -255
rect 401 -289 417 -255
rect 351 -323 417 -289
rect 351 -357 367 -323
rect 401 -357 417 -323
rect 351 -391 417 -357
rect 351 -425 367 -391
rect 401 -425 417 -391
rect 351 -459 417 -425
rect 351 -493 367 -459
rect 401 -493 417 -459
rect 351 -527 417 -493
rect 351 -561 367 -527
rect 401 -561 417 -527
rect 351 -595 417 -561
rect 351 -629 367 -595
rect 401 -629 417 -595
rect 351 -663 417 -629
rect 351 -697 367 -663
rect 401 -697 417 -663
rect 351 -731 417 -697
rect 351 -765 367 -731
rect 401 -765 417 -731
rect 351 -800 417 -765
rect 447 765 509 800
rect 447 731 463 765
rect 497 731 509 765
rect 447 697 509 731
rect 447 663 463 697
rect 497 663 509 697
rect 447 629 509 663
rect 447 595 463 629
rect 497 595 509 629
rect 447 561 509 595
rect 447 527 463 561
rect 497 527 509 561
rect 447 493 509 527
rect 447 459 463 493
rect 497 459 509 493
rect 447 425 509 459
rect 447 391 463 425
rect 497 391 509 425
rect 447 357 509 391
rect 447 323 463 357
rect 497 323 509 357
rect 447 289 509 323
rect 447 255 463 289
rect 497 255 509 289
rect 447 221 509 255
rect 447 187 463 221
rect 497 187 509 221
rect 447 153 509 187
rect 447 119 463 153
rect 497 119 509 153
rect 447 85 509 119
rect 447 51 463 85
rect 497 51 509 85
rect 447 17 509 51
rect 447 -17 463 17
rect 497 -17 509 17
rect 447 -51 509 -17
rect 447 -85 463 -51
rect 497 -85 509 -51
rect 447 -119 509 -85
rect 447 -153 463 -119
rect 497 -153 509 -119
rect 447 -187 509 -153
rect 447 -221 463 -187
rect 497 -221 509 -187
rect 447 -255 509 -221
rect 447 -289 463 -255
rect 497 -289 509 -255
rect 447 -323 509 -289
rect 447 -357 463 -323
rect 497 -357 509 -323
rect 447 -391 509 -357
rect 447 -425 463 -391
rect 497 -425 509 -391
rect 447 -459 509 -425
rect 447 -493 463 -459
rect 497 -493 509 -459
rect 447 -527 509 -493
rect 447 -561 463 -527
rect 497 -561 509 -527
rect 447 -595 509 -561
rect 447 -629 463 -595
rect 497 -629 509 -595
rect 447 -663 509 -629
rect 447 -697 463 -663
rect 497 -697 509 -663
rect 447 -731 509 -697
rect 447 -765 463 -731
rect 497 -765 509 -731
rect 447 -800 509 -765
<< pdiffc >>
rect -497 731 -463 765
rect -497 663 -463 697
rect -497 595 -463 629
rect -497 527 -463 561
rect -497 459 -463 493
rect -497 391 -463 425
rect -497 323 -463 357
rect -497 255 -463 289
rect -497 187 -463 221
rect -497 119 -463 153
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -497 -153 -463 -119
rect -497 -221 -463 -187
rect -497 -289 -463 -255
rect -497 -357 -463 -323
rect -497 -425 -463 -391
rect -497 -493 -463 -459
rect -497 -561 -463 -527
rect -497 -629 -463 -595
rect -497 -697 -463 -663
rect -497 -765 -463 -731
rect -401 731 -367 765
rect -401 663 -367 697
rect -401 595 -367 629
rect -401 527 -367 561
rect -401 459 -367 493
rect -401 391 -367 425
rect -401 323 -367 357
rect -401 255 -367 289
rect -401 187 -367 221
rect -401 119 -367 153
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -401 -153 -367 -119
rect -401 -221 -367 -187
rect -401 -289 -367 -255
rect -401 -357 -367 -323
rect -401 -425 -367 -391
rect -401 -493 -367 -459
rect -401 -561 -367 -527
rect -401 -629 -367 -595
rect -401 -697 -367 -663
rect -401 -765 -367 -731
rect -305 731 -271 765
rect -305 663 -271 697
rect -305 595 -271 629
rect -305 527 -271 561
rect -305 459 -271 493
rect -305 391 -271 425
rect -305 323 -271 357
rect -305 255 -271 289
rect -305 187 -271 221
rect -305 119 -271 153
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -305 -153 -271 -119
rect -305 -221 -271 -187
rect -305 -289 -271 -255
rect -305 -357 -271 -323
rect -305 -425 -271 -391
rect -305 -493 -271 -459
rect -305 -561 -271 -527
rect -305 -629 -271 -595
rect -305 -697 -271 -663
rect -305 -765 -271 -731
rect -209 731 -175 765
rect -209 663 -175 697
rect -209 595 -175 629
rect -209 527 -175 561
rect -209 459 -175 493
rect -209 391 -175 425
rect -209 323 -175 357
rect -209 255 -175 289
rect -209 187 -175 221
rect -209 119 -175 153
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -209 -153 -175 -119
rect -209 -221 -175 -187
rect -209 -289 -175 -255
rect -209 -357 -175 -323
rect -209 -425 -175 -391
rect -209 -493 -175 -459
rect -209 -561 -175 -527
rect -209 -629 -175 -595
rect -209 -697 -175 -663
rect -209 -765 -175 -731
rect -113 731 -79 765
rect -113 663 -79 697
rect -113 595 -79 629
rect -113 527 -79 561
rect -113 459 -79 493
rect -113 391 -79 425
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -113 -425 -79 -391
rect -113 -493 -79 -459
rect -113 -561 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -663
rect -113 -765 -79 -731
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect 79 731 113 765
rect 79 663 113 697
rect 79 595 113 629
rect 79 527 113 561
rect 79 459 113 493
rect 79 391 113 425
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 79 -425 113 -391
rect 79 -493 113 -459
rect 79 -561 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -663
rect 79 -765 113 -731
rect 175 731 209 765
rect 175 663 209 697
rect 175 595 209 629
rect 175 527 209 561
rect 175 459 209 493
rect 175 391 209 425
rect 175 323 209 357
rect 175 255 209 289
rect 175 187 209 221
rect 175 119 209 153
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 175 -153 209 -119
rect 175 -221 209 -187
rect 175 -289 209 -255
rect 175 -357 209 -323
rect 175 -425 209 -391
rect 175 -493 209 -459
rect 175 -561 209 -527
rect 175 -629 209 -595
rect 175 -697 209 -663
rect 175 -765 209 -731
rect 271 731 305 765
rect 271 663 305 697
rect 271 595 305 629
rect 271 527 305 561
rect 271 459 305 493
rect 271 391 305 425
rect 271 323 305 357
rect 271 255 305 289
rect 271 187 305 221
rect 271 119 305 153
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 271 -153 305 -119
rect 271 -221 305 -187
rect 271 -289 305 -255
rect 271 -357 305 -323
rect 271 -425 305 -391
rect 271 -493 305 -459
rect 271 -561 305 -527
rect 271 -629 305 -595
rect 271 -697 305 -663
rect 271 -765 305 -731
rect 367 731 401 765
rect 367 663 401 697
rect 367 595 401 629
rect 367 527 401 561
rect 367 459 401 493
rect 367 391 401 425
rect 367 323 401 357
rect 367 255 401 289
rect 367 187 401 221
rect 367 119 401 153
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 367 -153 401 -119
rect 367 -221 401 -187
rect 367 -289 401 -255
rect 367 -357 401 -323
rect 367 -425 401 -391
rect 367 -493 401 -459
rect 367 -561 401 -527
rect 367 -629 401 -595
rect 367 -697 401 -663
rect 367 -765 401 -731
rect 463 731 497 765
rect 463 663 497 697
rect 463 595 497 629
rect 463 527 497 561
rect 463 459 497 493
rect 463 391 497 425
rect 463 323 497 357
rect 463 255 497 289
rect 463 187 497 221
rect 463 119 497 153
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 463 -153 497 -119
rect 463 -221 497 -187
rect 463 -289 497 -255
rect 463 -357 497 -323
rect 463 -425 497 -391
rect 463 -493 497 -459
rect 463 -561 497 -527
rect 463 -629 497 -595
rect 463 -697 497 -663
rect 463 -765 497 -731
<< nsubdiff >>
rect -611 949 -493 983
rect -459 949 -425 983
rect -391 949 -357 983
rect -323 949 -289 983
rect -255 949 -221 983
rect -187 949 -153 983
rect -119 949 -85 983
rect -51 949 -17 983
rect 17 949 51 983
rect 85 949 119 983
rect 153 949 187 983
rect 221 949 255 983
rect 289 949 323 983
rect 357 949 391 983
rect 425 949 459 983
rect 493 949 611 983
rect -611 867 -577 949
rect -611 799 -577 833
rect 577 867 611 949
rect -611 731 -577 765
rect -611 663 -577 697
rect -611 595 -577 629
rect -611 527 -577 561
rect -611 459 -577 493
rect -611 391 -577 425
rect -611 323 -577 357
rect -611 255 -577 289
rect -611 187 -577 221
rect -611 119 -577 153
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect -611 -153 -577 -119
rect -611 -221 -577 -187
rect -611 -289 -577 -255
rect -611 -357 -577 -323
rect -611 -425 -577 -391
rect -611 -493 -577 -459
rect -611 -561 -577 -527
rect -611 -629 -577 -595
rect -611 -697 -577 -663
rect -611 -765 -577 -731
rect -611 -833 -577 -799
rect 577 799 611 833
rect 577 731 611 765
rect 577 663 611 697
rect 577 595 611 629
rect 577 527 611 561
rect 577 459 611 493
rect 577 391 611 425
rect 577 323 611 357
rect 577 255 611 289
rect 577 187 611 221
rect 577 119 611 153
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect 577 -153 611 -119
rect 577 -221 611 -187
rect 577 -289 611 -255
rect 577 -357 611 -323
rect 577 -425 611 -391
rect 577 -493 611 -459
rect 577 -561 611 -527
rect 577 -629 611 -595
rect 577 -697 611 -663
rect 577 -765 611 -731
rect -611 -949 -577 -867
rect 577 -833 611 -799
rect 577 -949 611 -867
rect -611 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 611 -949
<< nsubdiffcont >>
rect -493 949 -459 983
rect -425 949 -391 983
rect -357 949 -323 983
rect -289 949 -255 983
rect -221 949 -187 983
rect -153 949 -119 983
rect -85 949 -51 983
rect -17 949 17 983
rect 51 949 85 983
rect 119 949 153 983
rect 187 949 221 983
rect 255 949 289 983
rect 323 949 357 983
rect 391 949 425 983
rect 459 949 493 983
rect -611 833 -577 867
rect 577 833 611 867
rect -611 765 -577 799
rect -611 697 -577 731
rect -611 629 -577 663
rect -611 561 -577 595
rect -611 493 -577 527
rect -611 425 -577 459
rect -611 357 -577 391
rect -611 289 -577 323
rect -611 221 -577 255
rect -611 153 -577 187
rect -611 85 -577 119
rect -611 17 -577 51
rect -611 -51 -577 -17
rect -611 -119 -577 -85
rect -611 -187 -577 -153
rect -611 -255 -577 -221
rect -611 -323 -577 -289
rect -611 -391 -577 -357
rect -611 -459 -577 -425
rect -611 -527 -577 -493
rect -611 -595 -577 -561
rect -611 -663 -577 -629
rect -611 -731 -577 -697
rect -611 -799 -577 -765
rect 577 765 611 799
rect 577 697 611 731
rect 577 629 611 663
rect 577 561 611 595
rect 577 493 611 527
rect 577 425 611 459
rect 577 357 611 391
rect 577 289 611 323
rect 577 221 611 255
rect 577 153 611 187
rect 577 85 611 119
rect 577 17 611 51
rect 577 -51 611 -17
rect 577 -119 611 -85
rect 577 -187 611 -153
rect 577 -255 611 -221
rect 577 -323 611 -289
rect 577 -391 611 -357
rect 577 -459 611 -425
rect 577 -527 611 -493
rect 577 -595 611 -561
rect 577 -663 611 -629
rect 577 -731 611 -697
rect 577 -799 611 -765
rect -611 -867 -577 -833
rect 577 -867 611 -833
rect -493 -983 -459 -949
rect -425 -983 -391 -949
rect -357 -983 -323 -949
rect -289 -983 -255 -949
rect -221 -983 -187 -949
rect -153 -983 -119 -949
rect -85 -983 -51 -949
rect -17 -983 17 -949
rect 51 -983 85 -949
rect 119 -983 153 -949
rect 187 -983 221 -949
rect 255 -983 289 -949
rect 323 -983 357 -949
rect 391 -983 425 -949
rect 459 -983 493 -949
<< poly >>
rect -369 881 -303 897
rect -369 847 -353 881
rect -319 847 -303 881
rect -369 831 -303 847
rect -177 881 -111 897
rect -177 847 -161 881
rect -127 847 -111 881
rect -177 831 -111 847
rect 15 881 81 897
rect 15 847 31 881
rect 65 847 81 881
rect 15 831 81 847
rect 207 881 273 897
rect 207 847 223 881
rect 257 847 273 881
rect 207 831 273 847
rect 399 881 465 897
rect 399 847 415 881
rect 449 847 465 881
rect 399 831 465 847
rect -447 800 -417 826
rect -351 800 -321 831
rect -255 800 -225 826
rect -159 800 -129 831
rect -63 800 -33 826
rect 33 800 63 831
rect 129 800 159 826
rect 225 800 255 831
rect 321 800 351 826
rect 417 800 447 831
rect -447 -831 -417 -800
rect -351 -826 -321 -800
rect -255 -831 -225 -800
rect -159 -826 -129 -800
rect -63 -831 -33 -800
rect 33 -826 63 -800
rect 129 -831 159 -800
rect 225 -826 255 -800
rect 321 -831 351 -800
rect 417 -826 447 -800
rect -465 -847 -399 -831
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -465 -897 -399 -881
rect -273 -847 -207 -831
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -273 -897 -207 -881
rect -81 -847 -15 -831
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect -81 -897 -15 -881
rect 111 -847 177 -831
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 111 -897 177 -881
rect 303 -847 369 -831
rect 303 -881 319 -847
rect 353 -881 369 -847
rect 303 -897 369 -881
<< polycont >>
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
<< locali >>
rect -611 949 -493 983
rect -459 949 -425 983
rect -391 949 -357 983
rect -323 949 -289 983
rect -255 949 -221 983
rect -187 949 -153 983
rect -119 949 -85 983
rect -51 949 -17 983
rect 17 949 51 983
rect 85 949 119 983
rect 153 949 187 983
rect 221 949 255 983
rect 289 949 323 983
rect 357 949 391 983
rect 425 949 459 983
rect 493 949 611 983
rect -611 867 -577 949
rect -369 847 -353 881
rect -319 847 -303 881
rect -177 847 -161 881
rect -127 847 -111 881
rect 15 847 31 881
rect 65 847 81 881
rect 207 847 223 881
rect 257 847 273 881
rect 399 847 415 881
rect 449 847 465 881
rect 577 867 611 949
rect -611 799 -577 833
rect -611 731 -577 765
rect -611 663 -577 697
rect -611 595 -577 629
rect -611 527 -577 561
rect -611 459 -577 493
rect -611 391 -577 425
rect -611 323 -577 357
rect -611 255 -577 289
rect -611 187 -577 221
rect -611 119 -577 153
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect -611 -153 -577 -119
rect -611 -221 -577 -187
rect -611 -289 -577 -255
rect -611 -357 -577 -323
rect -611 -425 -577 -391
rect -611 -493 -577 -459
rect -611 -561 -577 -527
rect -611 -629 -577 -595
rect -611 -697 -577 -663
rect -611 -765 -577 -731
rect -611 -833 -577 -799
rect -497 773 -463 804
rect -497 701 -463 731
rect -497 629 -463 663
rect -497 561 -463 595
rect -497 493 -463 523
rect -497 425 -463 451
rect -497 357 -463 379
rect -497 289 -463 307
rect -497 221 -463 235
rect -497 153 -463 163
rect -497 85 -463 91
rect -497 17 -463 19
rect -497 -19 -463 -17
rect -497 -91 -463 -85
rect -497 -163 -463 -153
rect -497 -235 -463 -221
rect -497 -307 -463 -289
rect -497 -379 -463 -357
rect -497 -451 -463 -425
rect -497 -523 -463 -493
rect -497 -595 -463 -561
rect -497 -663 -463 -629
rect -497 -731 -463 -701
rect -497 -804 -463 -773
rect -401 773 -367 804
rect -401 701 -367 731
rect -401 629 -367 663
rect -401 561 -367 595
rect -401 493 -367 523
rect -401 425 -367 451
rect -401 357 -367 379
rect -401 289 -367 307
rect -401 221 -367 235
rect -401 153 -367 163
rect -401 85 -367 91
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -91 -367 -85
rect -401 -163 -367 -153
rect -401 -235 -367 -221
rect -401 -307 -367 -289
rect -401 -379 -367 -357
rect -401 -451 -367 -425
rect -401 -523 -367 -493
rect -401 -595 -367 -561
rect -401 -663 -367 -629
rect -401 -731 -367 -701
rect -401 -804 -367 -773
rect -305 773 -271 804
rect -305 701 -271 731
rect -305 629 -271 663
rect -305 561 -271 595
rect -305 493 -271 523
rect -305 425 -271 451
rect -305 357 -271 379
rect -305 289 -271 307
rect -305 221 -271 235
rect -305 153 -271 163
rect -305 85 -271 91
rect -305 17 -271 19
rect -305 -19 -271 -17
rect -305 -91 -271 -85
rect -305 -163 -271 -153
rect -305 -235 -271 -221
rect -305 -307 -271 -289
rect -305 -379 -271 -357
rect -305 -451 -271 -425
rect -305 -523 -271 -493
rect -305 -595 -271 -561
rect -305 -663 -271 -629
rect -305 -731 -271 -701
rect -305 -804 -271 -773
rect -209 773 -175 804
rect -209 701 -175 731
rect -209 629 -175 663
rect -209 561 -175 595
rect -209 493 -175 523
rect -209 425 -175 451
rect -209 357 -175 379
rect -209 289 -175 307
rect -209 221 -175 235
rect -209 153 -175 163
rect -209 85 -175 91
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -91 -175 -85
rect -209 -163 -175 -153
rect -209 -235 -175 -221
rect -209 -307 -175 -289
rect -209 -379 -175 -357
rect -209 -451 -175 -425
rect -209 -523 -175 -493
rect -209 -595 -175 -561
rect -209 -663 -175 -629
rect -209 -731 -175 -701
rect -209 -804 -175 -773
rect -113 773 -79 804
rect -113 701 -79 731
rect -113 629 -79 663
rect -113 561 -79 595
rect -113 493 -79 523
rect -113 425 -79 451
rect -113 357 -79 379
rect -113 289 -79 307
rect -113 221 -79 235
rect -113 153 -79 163
rect -113 85 -79 91
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -91 -79 -85
rect -113 -163 -79 -153
rect -113 -235 -79 -221
rect -113 -307 -79 -289
rect -113 -379 -79 -357
rect -113 -451 -79 -425
rect -113 -523 -79 -493
rect -113 -595 -79 -561
rect -113 -663 -79 -629
rect -113 -731 -79 -701
rect -113 -804 -79 -773
rect -17 773 17 804
rect -17 701 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -701
rect -17 -804 17 -773
rect 79 773 113 804
rect 79 701 113 731
rect 79 629 113 663
rect 79 561 113 595
rect 79 493 113 523
rect 79 425 113 451
rect 79 357 113 379
rect 79 289 113 307
rect 79 221 113 235
rect 79 153 113 163
rect 79 85 113 91
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -91 113 -85
rect 79 -163 113 -153
rect 79 -235 113 -221
rect 79 -307 113 -289
rect 79 -379 113 -357
rect 79 -451 113 -425
rect 79 -523 113 -493
rect 79 -595 113 -561
rect 79 -663 113 -629
rect 79 -731 113 -701
rect 79 -804 113 -773
rect 175 773 209 804
rect 175 701 209 731
rect 175 629 209 663
rect 175 561 209 595
rect 175 493 209 523
rect 175 425 209 451
rect 175 357 209 379
rect 175 289 209 307
rect 175 221 209 235
rect 175 153 209 163
rect 175 85 209 91
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -91 209 -85
rect 175 -163 209 -153
rect 175 -235 209 -221
rect 175 -307 209 -289
rect 175 -379 209 -357
rect 175 -451 209 -425
rect 175 -523 209 -493
rect 175 -595 209 -561
rect 175 -663 209 -629
rect 175 -731 209 -701
rect 175 -804 209 -773
rect 271 773 305 804
rect 271 701 305 731
rect 271 629 305 663
rect 271 561 305 595
rect 271 493 305 523
rect 271 425 305 451
rect 271 357 305 379
rect 271 289 305 307
rect 271 221 305 235
rect 271 153 305 163
rect 271 85 305 91
rect 271 17 305 19
rect 271 -19 305 -17
rect 271 -91 305 -85
rect 271 -163 305 -153
rect 271 -235 305 -221
rect 271 -307 305 -289
rect 271 -379 305 -357
rect 271 -451 305 -425
rect 271 -523 305 -493
rect 271 -595 305 -561
rect 271 -663 305 -629
rect 271 -731 305 -701
rect 271 -804 305 -773
rect 367 773 401 804
rect 367 701 401 731
rect 367 629 401 663
rect 367 561 401 595
rect 367 493 401 523
rect 367 425 401 451
rect 367 357 401 379
rect 367 289 401 307
rect 367 221 401 235
rect 367 153 401 163
rect 367 85 401 91
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -91 401 -85
rect 367 -163 401 -153
rect 367 -235 401 -221
rect 367 -307 401 -289
rect 367 -379 401 -357
rect 367 -451 401 -425
rect 367 -523 401 -493
rect 367 -595 401 -561
rect 367 -663 401 -629
rect 367 -731 401 -701
rect 367 -804 401 -773
rect 463 773 497 804
rect 463 701 497 731
rect 463 629 497 663
rect 463 561 497 595
rect 463 493 497 523
rect 463 425 497 451
rect 463 357 497 379
rect 463 289 497 307
rect 463 221 497 235
rect 463 153 497 163
rect 463 85 497 91
rect 463 17 497 19
rect 463 -19 497 -17
rect 463 -91 497 -85
rect 463 -163 497 -153
rect 463 -235 497 -221
rect 463 -307 497 -289
rect 463 -379 497 -357
rect 463 -451 497 -425
rect 463 -523 497 -493
rect 463 -595 497 -561
rect 463 -663 497 -629
rect 463 -731 497 -701
rect 463 -804 497 -773
rect 577 799 611 833
rect 577 731 611 765
rect 577 663 611 697
rect 577 595 611 629
rect 577 527 611 561
rect 577 459 611 493
rect 577 391 611 425
rect 577 323 611 357
rect 577 255 611 289
rect 577 187 611 221
rect 577 119 611 153
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect 577 -153 611 -119
rect 577 -221 611 -187
rect 577 -289 611 -255
rect 577 -357 611 -323
rect 577 -425 611 -391
rect 577 -493 611 -459
rect 577 -561 611 -527
rect 577 -629 611 -595
rect 577 -697 611 -663
rect 577 -765 611 -731
rect 577 -833 611 -799
rect -611 -949 -577 -867
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 303 -881 319 -847
rect 353 -881 369 -847
rect 577 -949 611 -867
rect -611 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 611 -949
<< viali >>
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect -497 765 -463 773
rect -497 739 -463 765
rect -497 697 -463 701
rect -497 667 -463 697
rect -497 595 -463 629
rect -497 527 -463 557
rect -497 523 -463 527
rect -497 459 -463 485
rect -497 451 -463 459
rect -497 391 -463 413
rect -497 379 -463 391
rect -497 323 -463 341
rect -497 307 -463 323
rect -497 255 -463 269
rect -497 235 -463 255
rect -497 187 -463 197
rect -497 163 -463 187
rect -497 119 -463 125
rect -497 91 -463 119
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -497 -119 -463 -91
rect -497 -125 -463 -119
rect -497 -187 -463 -163
rect -497 -197 -463 -187
rect -497 -255 -463 -235
rect -497 -269 -463 -255
rect -497 -323 -463 -307
rect -497 -341 -463 -323
rect -497 -391 -463 -379
rect -497 -413 -463 -391
rect -497 -459 -463 -451
rect -497 -485 -463 -459
rect -497 -527 -463 -523
rect -497 -557 -463 -527
rect -497 -629 -463 -595
rect -497 -697 -463 -667
rect -497 -701 -463 -697
rect -497 -765 -463 -739
rect -497 -773 -463 -765
rect -401 765 -367 773
rect -401 739 -367 765
rect -401 697 -367 701
rect -401 667 -367 697
rect -401 595 -367 629
rect -401 527 -367 557
rect -401 523 -367 527
rect -401 459 -367 485
rect -401 451 -367 459
rect -401 391 -367 413
rect -401 379 -367 391
rect -401 323 -367 341
rect -401 307 -367 323
rect -401 255 -367 269
rect -401 235 -367 255
rect -401 187 -367 197
rect -401 163 -367 187
rect -401 119 -367 125
rect -401 91 -367 119
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -401 -119 -367 -91
rect -401 -125 -367 -119
rect -401 -187 -367 -163
rect -401 -197 -367 -187
rect -401 -255 -367 -235
rect -401 -269 -367 -255
rect -401 -323 -367 -307
rect -401 -341 -367 -323
rect -401 -391 -367 -379
rect -401 -413 -367 -391
rect -401 -459 -367 -451
rect -401 -485 -367 -459
rect -401 -527 -367 -523
rect -401 -557 -367 -527
rect -401 -629 -367 -595
rect -401 -697 -367 -667
rect -401 -701 -367 -697
rect -401 -765 -367 -739
rect -401 -773 -367 -765
rect -305 765 -271 773
rect -305 739 -271 765
rect -305 697 -271 701
rect -305 667 -271 697
rect -305 595 -271 629
rect -305 527 -271 557
rect -305 523 -271 527
rect -305 459 -271 485
rect -305 451 -271 459
rect -305 391 -271 413
rect -305 379 -271 391
rect -305 323 -271 341
rect -305 307 -271 323
rect -305 255 -271 269
rect -305 235 -271 255
rect -305 187 -271 197
rect -305 163 -271 187
rect -305 119 -271 125
rect -305 91 -271 119
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -305 -119 -271 -91
rect -305 -125 -271 -119
rect -305 -187 -271 -163
rect -305 -197 -271 -187
rect -305 -255 -271 -235
rect -305 -269 -271 -255
rect -305 -323 -271 -307
rect -305 -341 -271 -323
rect -305 -391 -271 -379
rect -305 -413 -271 -391
rect -305 -459 -271 -451
rect -305 -485 -271 -459
rect -305 -527 -271 -523
rect -305 -557 -271 -527
rect -305 -629 -271 -595
rect -305 -697 -271 -667
rect -305 -701 -271 -697
rect -305 -765 -271 -739
rect -305 -773 -271 -765
rect -209 765 -175 773
rect -209 739 -175 765
rect -209 697 -175 701
rect -209 667 -175 697
rect -209 595 -175 629
rect -209 527 -175 557
rect -209 523 -175 527
rect -209 459 -175 485
rect -209 451 -175 459
rect -209 391 -175 413
rect -209 379 -175 391
rect -209 323 -175 341
rect -209 307 -175 323
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -209 -323 -175 -307
rect -209 -341 -175 -323
rect -209 -391 -175 -379
rect -209 -413 -175 -391
rect -209 -459 -175 -451
rect -209 -485 -175 -459
rect -209 -527 -175 -523
rect -209 -557 -175 -527
rect -209 -629 -175 -595
rect -209 -697 -175 -667
rect -209 -701 -175 -697
rect -209 -765 -175 -739
rect -209 -773 -175 -765
rect -113 765 -79 773
rect -113 739 -79 765
rect -113 697 -79 701
rect -113 667 -79 697
rect -113 595 -79 629
rect -113 527 -79 557
rect -113 523 -79 527
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -113 -527 -79 -523
rect -113 -557 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -667
rect -113 -701 -79 -697
rect -113 -765 -79 -739
rect -113 -773 -79 -765
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect 79 765 113 773
rect 79 739 113 765
rect 79 697 113 701
rect 79 667 113 697
rect 79 595 113 629
rect 79 527 113 557
rect 79 523 113 527
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 79 -527 113 -523
rect 79 -557 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -667
rect 79 -701 113 -697
rect 79 -765 113 -739
rect 79 -773 113 -765
rect 175 765 209 773
rect 175 739 209 765
rect 175 697 209 701
rect 175 667 209 697
rect 175 595 209 629
rect 175 527 209 557
rect 175 523 209 527
rect 175 459 209 485
rect 175 451 209 459
rect 175 391 209 413
rect 175 379 209 391
rect 175 323 209 341
rect 175 307 209 323
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect 175 -323 209 -307
rect 175 -341 209 -323
rect 175 -391 209 -379
rect 175 -413 209 -391
rect 175 -459 209 -451
rect 175 -485 209 -459
rect 175 -527 209 -523
rect 175 -557 209 -527
rect 175 -629 209 -595
rect 175 -697 209 -667
rect 175 -701 209 -697
rect 175 -765 209 -739
rect 175 -773 209 -765
rect 271 765 305 773
rect 271 739 305 765
rect 271 697 305 701
rect 271 667 305 697
rect 271 595 305 629
rect 271 527 305 557
rect 271 523 305 527
rect 271 459 305 485
rect 271 451 305 459
rect 271 391 305 413
rect 271 379 305 391
rect 271 323 305 341
rect 271 307 305 323
rect 271 255 305 269
rect 271 235 305 255
rect 271 187 305 197
rect 271 163 305 187
rect 271 119 305 125
rect 271 91 305 119
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 271 -119 305 -91
rect 271 -125 305 -119
rect 271 -187 305 -163
rect 271 -197 305 -187
rect 271 -255 305 -235
rect 271 -269 305 -255
rect 271 -323 305 -307
rect 271 -341 305 -323
rect 271 -391 305 -379
rect 271 -413 305 -391
rect 271 -459 305 -451
rect 271 -485 305 -459
rect 271 -527 305 -523
rect 271 -557 305 -527
rect 271 -629 305 -595
rect 271 -697 305 -667
rect 271 -701 305 -697
rect 271 -765 305 -739
rect 271 -773 305 -765
rect 367 765 401 773
rect 367 739 401 765
rect 367 697 401 701
rect 367 667 401 697
rect 367 595 401 629
rect 367 527 401 557
rect 367 523 401 527
rect 367 459 401 485
rect 367 451 401 459
rect 367 391 401 413
rect 367 379 401 391
rect 367 323 401 341
rect 367 307 401 323
rect 367 255 401 269
rect 367 235 401 255
rect 367 187 401 197
rect 367 163 401 187
rect 367 119 401 125
rect 367 91 401 119
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 367 -119 401 -91
rect 367 -125 401 -119
rect 367 -187 401 -163
rect 367 -197 401 -187
rect 367 -255 401 -235
rect 367 -269 401 -255
rect 367 -323 401 -307
rect 367 -341 401 -323
rect 367 -391 401 -379
rect 367 -413 401 -391
rect 367 -459 401 -451
rect 367 -485 401 -459
rect 367 -527 401 -523
rect 367 -557 401 -527
rect 367 -629 401 -595
rect 367 -697 401 -667
rect 367 -701 401 -697
rect 367 -765 401 -739
rect 367 -773 401 -765
rect 463 765 497 773
rect 463 739 497 765
rect 463 697 497 701
rect 463 667 497 697
rect 463 595 497 629
rect 463 527 497 557
rect 463 523 497 527
rect 463 459 497 485
rect 463 451 497 459
rect 463 391 497 413
rect 463 379 497 391
rect 463 323 497 341
rect 463 307 497 323
rect 463 255 497 269
rect 463 235 497 255
rect 463 187 497 197
rect 463 163 497 187
rect 463 119 497 125
rect 463 91 497 119
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 463 -119 497 -91
rect 463 -125 497 -119
rect 463 -187 497 -163
rect 463 -197 497 -187
rect 463 -255 497 -235
rect 463 -269 497 -255
rect 463 -323 497 -307
rect 463 -341 497 -323
rect 463 -391 497 -379
rect 463 -413 497 -391
rect 463 -459 497 -451
rect 463 -485 497 -459
rect 463 -527 497 -523
rect 463 -557 497 -527
rect 463 -629 497 -595
rect 463 -697 497 -667
rect 463 -701 497 -697
rect 463 -765 497 -739
rect 463 -773 497 -765
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
<< metal1 >>
rect -365 881 -307 887
rect -365 847 -353 881
rect -319 847 -307 881
rect -365 841 -307 847
rect -173 881 -115 887
rect -173 847 -161 881
rect -127 847 -115 881
rect -173 841 -115 847
rect 19 881 77 887
rect 19 847 31 881
rect 65 847 77 881
rect 19 841 77 847
rect 211 881 269 887
rect 211 847 223 881
rect 257 847 269 881
rect 211 841 269 847
rect 403 881 461 887
rect 403 847 415 881
rect 449 847 461 881
rect 403 841 461 847
rect -503 773 -457 800
rect -503 739 -497 773
rect -463 739 -457 773
rect -503 701 -457 739
rect -503 667 -497 701
rect -463 667 -457 701
rect -503 629 -457 667
rect -503 595 -497 629
rect -463 595 -457 629
rect -503 557 -457 595
rect -503 523 -497 557
rect -463 523 -457 557
rect -503 485 -457 523
rect -503 451 -497 485
rect -463 451 -457 485
rect -503 413 -457 451
rect -503 379 -497 413
rect -463 379 -457 413
rect -503 341 -457 379
rect -503 307 -497 341
rect -463 307 -457 341
rect -503 269 -457 307
rect -503 235 -497 269
rect -463 235 -457 269
rect -503 197 -457 235
rect -503 163 -497 197
rect -463 163 -457 197
rect -503 125 -457 163
rect -503 91 -497 125
rect -463 91 -457 125
rect -503 53 -457 91
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -91 -457 -53
rect -503 -125 -497 -91
rect -463 -125 -457 -91
rect -503 -163 -457 -125
rect -503 -197 -497 -163
rect -463 -197 -457 -163
rect -503 -235 -457 -197
rect -503 -269 -497 -235
rect -463 -269 -457 -235
rect -503 -307 -457 -269
rect -503 -341 -497 -307
rect -463 -341 -457 -307
rect -503 -379 -457 -341
rect -503 -413 -497 -379
rect -463 -413 -457 -379
rect -503 -451 -457 -413
rect -503 -485 -497 -451
rect -463 -485 -457 -451
rect -503 -523 -457 -485
rect -503 -557 -497 -523
rect -463 -557 -457 -523
rect -503 -595 -457 -557
rect -503 -629 -497 -595
rect -463 -629 -457 -595
rect -503 -667 -457 -629
rect -503 -701 -497 -667
rect -463 -701 -457 -667
rect -503 -739 -457 -701
rect -503 -773 -497 -739
rect -463 -773 -457 -739
rect -503 -800 -457 -773
rect -407 773 -361 800
rect -407 739 -401 773
rect -367 739 -361 773
rect -407 701 -361 739
rect -407 667 -401 701
rect -367 667 -361 701
rect -407 629 -361 667
rect -407 595 -401 629
rect -367 595 -361 629
rect -407 557 -361 595
rect -407 523 -401 557
rect -367 523 -361 557
rect -407 485 -361 523
rect -407 451 -401 485
rect -367 451 -361 485
rect -407 413 -361 451
rect -407 379 -401 413
rect -367 379 -361 413
rect -407 341 -361 379
rect -407 307 -401 341
rect -367 307 -361 341
rect -407 269 -361 307
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -307 -361 -269
rect -407 -341 -401 -307
rect -367 -341 -361 -307
rect -407 -379 -361 -341
rect -407 -413 -401 -379
rect -367 -413 -361 -379
rect -407 -451 -361 -413
rect -407 -485 -401 -451
rect -367 -485 -361 -451
rect -407 -523 -361 -485
rect -407 -557 -401 -523
rect -367 -557 -361 -523
rect -407 -595 -361 -557
rect -407 -629 -401 -595
rect -367 -629 -361 -595
rect -407 -667 -361 -629
rect -407 -701 -401 -667
rect -367 -701 -361 -667
rect -407 -739 -361 -701
rect -407 -773 -401 -739
rect -367 -773 -361 -739
rect -407 -800 -361 -773
rect -311 773 -265 800
rect -311 739 -305 773
rect -271 739 -265 773
rect -311 701 -265 739
rect -311 667 -305 701
rect -271 667 -265 701
rect -311 629 -265 667
rect -311 595 -305 629
rect -271 595 -265 629
rect -311 557 -265 595
rect -311 523 -305 557
rect -271 523 -265 557
rect -311 485 -265 523
rect -311 451 -305 485
rect -271 451 -265 485
rect -311 413 -265 451
rect -311 379 -305 413
rect -271 379 -265 413
rect -311 341 -265 379
rect -311 307 -305 341
rect -271 307 -265 341
rect -311 269 -265 307
rect -311 235 -305 269
rect -271 235 -265 269
rect -311 197 -265 235
rect -311 163 -305 197
rect -271 163 -265 197
rect -311 125 -265 163
rect -311 91 -305 125
rect -271 91 -265 125
rect -311 53 -265 91
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -91 -265 -53
rect -311 -125 -305 -91
rect -271 -125 -265 -91
rect -311 -163 -265 -125
rect -311 -197 -305 -163
rect -271 -197 -265 -163
rect -311 -235 -265 -197
rect -311 -269 -305 -235
rect -271 -269 -265 -235
rect -311 -307 -265 -269
rect -311 -341 -305 -307
rect -271 -341 -265 -307
rect -311 -379 -265 -341
rect -311 -413 -305 -379
rect -271 -413 -265 -379
rect -311 -451 -265 -413
rect -311 -485 -305 -451
rect -271 -485 -265 -451
rect -311 -523 -265 -485
rect -311 -557 -305 -523
rect -271 -557 -265 -523
rect -311 -595 -265 -557
rect -311 -629 -305 -595
rect -271 -629 -265 -595
rect -311 -667 -265 -629
rect -311 -701 -305 -667
rect -271 -701 -265 -667
rect -311 -739 -265 -701
rect -311 -773 -305 -739
rect -271 -773 -265 -739
rect -311 -800 -265 -773
rect -215 773 -169 800
rect -215 739 -209 773
rect -175 739 -169 773
rect -215 701 -169 739
rect -215 667 -209 701
rect -175 667 -169 701
rect -215 629 -169 667
rect -215 595 -209 629
rect -175 595 -169 629
rect -215 557 -169 595
rect -215 523 -209 557
rect -175 523 -169 557
rect -215 485 -169 523
rect -215 451 -209 485
rect -175 451 -169 485
rect -215 413 -169 451
rect -215 379 -209 413
rect -175 379 -169 413
rect -215 341 -169 379
rect -215 307 -209 341
rect -175 307 -169 341
rect -215 269 -169 307
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -307 -169 -269
rect -215 -341 -209 -307
rect -175 -341 -169 -307
rect -215 -379 -169 -341
rect -215 -413 -209 -379
rect -175 -413 -169 -379
rect -215 -451 -169 -413
rect -215 -485 -209 -451
rect -175 -485 -169 -451
rect -215 -523 -169 -485
rect -215 -557 -209 -523
rect -175 -557 -169 -523
rect -215 -595 -169 -557
rect -215 -629 -209 -595
rect -175 -629 -169 -595
rect -215 -667 -169 -629
rect -215 -701 -209 -667
rect -175 -701 -169 -667
rect -215 -739 -169 -701
rect -215 -773 -209 -739
rect -175 -773 -169 -739
rect -215 -800 -169 -773
rect -119 773 -73 800
rect -119 739 -113 773
rect -79 739 -73 773
rect -119 701 -73 739
rect -119 667 -113 701
rect -79 667 -73 701
rect -119 629 -73 667
rect -119 595 -113 629
rect -79 595 -73 629
rect -119 557 -73 595
rect -119 523 -113 557
rect -79 523 -73 557
rect -119 485 -73 523
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -523 -73 -485
rect -119 -557 -113 -523
rect -79 -557 -73 -523
rect -119 -595 -73 -557
rect -119 -629 -113 -595
rect -79 -629 -73 -595
rect -119 -667 -73 -629
rect -119 -701 -113 -667
rect -79 -701 -73 -667
rect -119 -739 -73 -701
rect -119 -773 -113 -739
rect -79 -773 -73 -739
rect -119 -800 -73 -773
rect -23 773 23 800
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -800 23 -773
rect 73 773 119 800
rect 73 739 79 773
rect 113 739 119 773
rect 73 701 119 739
rect 73 667 79 701
rect 113 667 119 701
rect 73 629 119 667
rect 73 595 79 629
rect 113 595 119 629
rect 73 557 119 595
rect 73 523 79 557
rect 113 523 119 557
rect 73 485 119 523
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -523 119 -485
rect 73 -557 79 -523
rect 113 -557 119 -523
rect 73 -595 119 -557
rect 73 -629 79 -595
rect 113 -629 119 -595
rect 73 -667 119 -629
rect 73 -701 79 -667
rect 113 -701 119 -667
rect 73 -739 119 -701
rect 73 -773 79 -739
rect 113 -773 119 -739
rect 73 -800 119 -773
rect 169 773 215 800
rect 169 739 175 773
rect 209 739 215 773
rect 169 701 215 739
rect 169 667 175 701
rect 209 667 215 701
rect 169 629 215 667
rect 169 595 175 629
rect 209 595 215 629
rect 169 557 215 595
rect 169 523 175 557
rect 209 523 215 557
rect 169 485 215 523
rect 169 451 175 485
rect 209 451 215 485
rect 169 413 215 451
rect 169 379 175 413
rect 209 379 215 413
rect 169 341 215 379
rect 169 307 175 341
rect 209 307 215 341
rect 169 269 215 307
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -307 215 -269
rect 169 -341 175 -307
rect 209 -341 215 -307
rect 169 -379 215 -341
rect 169 -413 175 -379
rect 209 -413 215 -379
rect 169 -451 215 -413
rect 169 -485 175 -451
rect 209 -485 215 -451
rect 169 -523 215 -485
rect 169 -557 175 -523
rect 209 -557 215 -523
rect 169 -595 215 -557
rect 169 -629 175 -595
rect 209 -629 215 -595
rect 169 -667 215 -629
rect 169 -701 175 -667
rect 209 -701 215 -667
rect 169 -739 215 -701
rect 169 -773 175 -739
rect 209 -773 215 -739
rect 169 -800 215 -773
rect 265 773 311 800
rect 265 739 271 773
rect 305 739 311 773
rect 265 701 311 739
rect 265 667 271 701
rect 305 667 311 701
rect 265 629 311 667
rect 265 595 271 629
rect 305 595 311 629
rect 265 557 311 595
rect 265 523 271 557
rect 305 523 311 557
rect 265 485 311 523
rect 265 451 271 485
rect 305 451 311 485
rect 265 413 311 451
rect 265 379 271 413
rect 305 379 311 413
rect 265 341 311 379
rect 265 307 271 341
rect 305 307 311 341
rect 265 269 311 307
rect 265 235 271 269
rect 305 235 311 269
rect 265 197 311 235
rect 265 163 271 197
rect 305 163 311 197
rect 265 125 311 163
rect 265 91 271 125
rect 305 91 311 125
rect 265 53 311 91
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -91 311 -53
rect 265 -125 271 -91
rect 305 -125 311 -91
rect 265 -163 311 -125
rect 265 -197 271 -163
rect 305 -197 311 -163
rect 265 -235 311 -197
rect 265 -269 271 -235
rect 305 -269 311 -235
rect 265 -307 311 -269
rect 265 -341 271 -307
rect 305 -341 311 -307
rect 265 -379 311 -341
rect 265 -413 271 -379
rect 305 -413 311 -379
rect 265 -451 311 -413
rect 265 -485 271 -451
rect 305 -485 311 -451
rect 265 -523 311 -485
rect 265 -557 271 -523
rect 305 -557 311 -523
rect 265 -595 311 -557
rect 265 -629 271 -595
rect 305 -629 311 -595
rect 265 -667 311 -629
rect 265 -701 271 -667
rect 305 -701 311 -667
rect 265 -739 311 -701
rect 265 -773 271 -739
rect 305 -773 311 -739
rect 265 -800 311 -773
rect 361 773 407 800
rect 361 739 367 773
rect 401 739 407 773
rect 361 701 407 739
rect 361 667 367 701
rect 401 667 407 701
rect 361 629 407 667
rect 361 595 367 629
rect 401 595 407 629
rect 361 557 407 595
rect 361 523 367 557
rect 401 523 407 557
rect 361 485 407 523
rect 361 451 367 485
rect 401 451 407 485
rect 361 413 407 451
rect 361 379 367 413
rect 401 379 407 413
rect 361 341 407 379
rect 361 307 367 341
rect 401 307 407 341
rect 361 269 407 307
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -307 407 -269
rect 361 -341 367 -307
rect 401 -341 407 -307
rect 361 -379 407 -341
rect 361 -413 367 -379
rect 401 -413 407 -379
rect 361 -451 407 -413
rect 361 -485 367 -451
rect 401 -485 407 -451
rect 361 -523 407 -485
rect 361 -557 367 -523
rect 401 -557 407 -523
rect 361 -595 407 -557
rect 361 -629 367 -595
rect 401 -629 407 -595
rect 361 -667 407 -629
rect 361 -701 367 -667
rect 401 -701 407 -667
rect 361 -739 407 -701
rect 361 -773 367 -739
rect 401 -773 407 -739
rect 361 -800 407 -773
rect 457 773 503 800
rect 457 739 463 773
rect 497 739 503 773
rect 457 701 503 739
rect 457 667 463 701
rect 497 667 503 701
rect 457 629 503 667
rect 457 595 463 629
rect 497 595 503 629
rect 457 557 503 595
rect 457 523 463 557
rect 497 523 503 557
rect 457 485 503 523
rect 457 451 463 485
rect 497 451 503 485
rect 457 413 503 451
rect 457 379 463 413
rect 497 379 503 413
rect 457 341 503 379
rect 457 307 463 341
rect 497 307 503 341
rect 457 269 503 307
rect 457 235 463 269
rect 497 235 503 269
rect 457 197 503 235
rect 457 163 463 197
rect 497 163 503 197
rect 457 125 503 163
rect 457 91 463 125
rect 497 91 503 125
rect 457 53 503 91
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -91 503 -53
rect 457 -125 463 -91
rect 497 -125 503 -91
rect 457 -163 503 -125
rect 457 -197 463 -163
rect 497 -197 503 -163
rect 457 -235 503 -197
rect 457 -269 463 -235
rect 497 -269 503 -235
rect 457 -307 503 -269
rect 457 -341 463 -307
rect 497 -341 503 -307
rect 457 -379 503 -341
rect 457 -413 463 -379
rect 497 -413 503 -379
rect 457 -451 503 -413
rect 457 -485 463 -451
rect 497 -485 503 -451
rect 457 -523 503 -485
rect 457 -557 463 -523
rect 497 -557 503 -523
rect 457 -595 503 -557
rect 457 -629 463 -595
rect 497 -629 503 -595
rect 457 -667 503 -629
rect 457 -701 463 -667
rect 497 -701 503 -667
rect 457 -739 503 -701
rect 457 -773 463 -739
rect 497 -773 503 -739
rect 457 -800 503 -773
rect -461 -847 -403 -841
rect -461 -881 -449 -847
rect -415 -881 -403 -847
rect -461 -887 -403 -881
rect -269 -847 -211 -841
rect -269 -881 -257 -847
rect -223 -881 -211 -847
rect -269 -887 -211 -881
rect -77 -847 -19 -841
rect -77 -881 -65 -847
rect -31 -881 -19 -847
rect -77 -887 -19 -881
rect 115 -847 173 -841
rect 115 -881 127 -847
rect 161 -881 173 -847
rect 115 -887 173 -881
rect 307 -847 365 -841
rect 307 -881 319 -847
rect 353 -881 365 -847
rect 307 -887 365 -881
<< properties >>
string FIXED_BBOX -594 -966 594 966
<< end >>
