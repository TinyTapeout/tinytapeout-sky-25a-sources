// Generated from: 20250609-161054_binTestAcc9611_seed571850_epochs50_2x1280_b256_lr75_interconnect.pth

module net (
    input  wire [255:0] in,
    output wire [1279:0] out,
    output wire [1269:0] categories
);
    wire [1280:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = ~(in[74] & in[165]); 
    assign layer_0[1] = in[138] & ~in[107]; 
    assign layer_0[2] = ~(in[135] | in[196]); 
    assign layer_0[3] = in[42] | in[197]; 
    assign layer_0[4] = in[75] & ~in[106]; 
    assign layer_0[5] = in[203] ^ in[154]; 
    assign layer_0[6] = in[159] ^ in[196]; 
    assign layer_0[7] = in[51] ^ in[40]; 
    assign layer_0[8] = ~(in[115] | in[116]); 
    assign layer_0[9] = in[149] & in[165]; 
    assign layer_0[10] = ~(in[156] | in[246]); 
    assign layer_0[11] = in[195] ^ in[133]; 
    assign layer_0[12] = in[202] ^ in[157]; 
    assign layer_0[13] = in[82] ^ in[51]; 
    assign layer_0[14] = in[103] ^ in[117]; 
    assign layer_0[15] = in[68]; 
    assign layer_0[16] = in[171] ^ in[194]; 
    assign layer_0[17] = in[124] ^ in[93]; 
    assign layer_0[18] = in[181]; 
    assign layer_0[19] = ~(in[87] ^ in[181]); 
    assign layer_0[20] = in[87] ^ in[39]; 
    assign layer_0[21] = ~in[155] | (in[220] & in[155]); 
    assign layer_0[22] = ~(in[91] | in[93]); 
    assign layer_0[23] = in[107] & ~in[122]; 
    assign layer_0[24] = in[40] & ~in[75]; 
    assign layer_0[25] = in[171] ^ in[218]; 
    assign layer_0[26] = in[89] | in[91]; 
    assign layer_0[27] = in[148] ^ in[127]; 
    assign layer_0[28] = ~(in[246] ^ in[172]); 
    assign layer_0[29] = ~(in[118] | in[116]); 
    assign layer_0[30] = in[230] | in[227]; 
    assign layer_0[31] = ~(in[26] | in[29]); 
    assign layer_0[32] = in[202] ^ in[228]; 
    assign layer_0[33] = ~(in[188] ^ in[155]); 
    assign layer_0[34] = in[70] & ~in[173]; 
    assign layer_0[35] = ~(in[88] ^ in[90]); 
    assign layer_0[36] = ~(in[84] ^ in[53]); 
    assign layer_0[37] = in[62] | in[185]; 
    assign layer_0[38] = ~(in[171] & in[140]); 
    assign layer_0[39] = in[219]; 
    assign layer_0[40] = ~(in[204] ^ in[202]); 
    assign layer_0[41] = in[51] | in[107]; 
    assign layer_0[42] = ~(in[133] | in[246]); 
    assign layer_0[43] = ~(in[71] ^ in[188]); 
    assign layer_0[44] = in[198] ^ in[188]; 
    assign layer_0[45] = ~(in[195] | in[213]); 
    assign layer_0[46] = ~(in[118] | in[95]); 
    assign layer_0[47] = in[134] | in[124]; 
    assign layer_0[48] = ~(in[91] | in[251]); 
    assign layer_0[49] = in[198] | in[125]; 
    assign layer_0[50] = ~(in[249] | in[82]); 
    assign layer_0[51] = in[54] ^ in[85]; 
    assign layer_0[52] = in[37] ^ in[68]; 
    assign layer_0[53] = in[147] ^ in[41]; 
    assign layer_0[54] = ~in[182]; 
    assign layer_0[55] = ~(in[24] ^ in[82]); 
    assign layer_0[56] = ~(in[203] | in[230]); 
    assign layer_0[57] = ~(in[155] & in[138]); 
    assign layer_0[58] = in[166] & ~in[88]; 
    assign layer_0[59] = in[180] | in[217]; 
    assign layer_0[60] = in[152] | in[121]; 
    assign layer_0[61] = ~(in[131] ^ in[118]); 
    assign layer_0[62] = ~in[119]; 
    assign layer_0[63] = ~(in[156] | in[139]); 
    assign layer_0[64] = ~in[185] | (in[139] & in[185]); 
    assign layer_0[65] = ~in[213] | (in[54] & in[213]); 
    assign layer_0[66] = in[125]; 
    assign layer_0[67] = ~in[198]; 
    assign layer_0[68] = in[206] ^ in[100]; 
    assign layer_0[69] = ~(in[178] ^ in[125]); 
    assign layer_0[70] = ~(in[125] ^ in[28]); 
    assign layer_0[71] = in[216] & in[154]; 
    assign layer_0[72] = ~(in[40] | in[84]); 
    assign layer_0[73] = in[132] & ~in[199]; 
    assign layer_0[74] = ~(in[187] ^ in[196]); 
    assign layer_0[75] = ~(in[218] ^ in[199]); 
    assign layer_0[76] = in[170] ^ in[172]; 
    assign layer_0[77] = ~(in[162] ^ in[249]); 
    assign layer_0[78] = ~in[38]; 
    assign layer_0[79] = ~(in[20] | in[181]); 
    assign layer_0[80] = ~(in[75] | in[58]); 
    assign layer_0[81] = in[119] ^ in[168]; 
    assign layer_0[82] = ~in[132] | (in[118] & in[132]); 
    assign layer_0[83] = in[60] ^ in[93]; 
    assign layer_0[84] = ~(in[106] ^ in[74]); 
    assign layer_0[85] = in[185]; 
    assign layer_0[86] = in[165] & ~in[155]; 
    assign layer_0[87] = ~(in[44] ^ in[73]); 
    assign layer_0[88] = in[28] ^ in[45]; 
    assign layer_0[89] = in[73] & ~in[212]; 
    assign layer_0[90] = in[73] & ~in[188]; 
    assign layer_0[91] = ~(in[228] | in[178]); 
    assign layer_0[92] = ~(in[190] ^ in[103]); 
    assign layer_0[93] = ~(in[38] | in[23]); 
    assign layer_0[94] = ~in[148]; 
    assign layer_0[95] = in[199] | in[214]; 
    assign layer_0[96] = ~(in[124] | in[78]); 
    assign layer_0[97] = in[69] | in[55]; 
    assign layer_0[98] = in[58] ^ in[54]; 
    assign layer_0[99] = in[102] ^ in[115]; 
    assign layer_0[100] = ~(in[138] | in[138]); 
    assign layer_0[101] = ~(in[106] | in[105]); 
    assign layer_0[102] = in[102] | in[100]; 
    assign layer_0[103] = in[150] ^ in[68]; 
    assign layer_0[104] = ~(in[118] ^ in[101]); 
    assign layer_0[105] = ~(in[156] | in[172]); 
    assign layer_0[106] = ~in[181] | (in[181] & in[227]); 
    assign layer_0[107] = in[212] & in[68]; 
    assign layer_0[108] = ~(in[139] ^ in[107]); 
    assign layer_0[109] = ~(in[21] | in[99]); 
    assign layer_0[110] = ~(in[163] | in[165]); 
    assign layer_0[111] = in[22] | in[221]; 
    assign layer_0[112] = in[54] & ~in[123]; 
    assign layer_0[113] = ~(in[124] | in[114]); 
    assign layer_0[114] = in[215] & ~in[153]; 
    assign layer_0[115] = in[148] & ~in[166]; 
    assign layer_0[116] = ~in[149]; 
    assign layer_0[117] = in[103] & ~in[248]; 
    assign layer_0[118] = in[56] & ~in[125]; 
    assign layer_0[119] = ~(in[196] ^ in[39]); 
    assign layer_0[120] = ~(in[121] ^ in[140]); 
    assign layer_0[121] = in[136] ^ in[84]; 
    assign layer_0[122] = ~(in[126] ^ in[108]); 
    assign layer_0[123] = ~(in[164] | in[167]); 
    assign layer_0[124] = in[171] ^ in[218]; 
    assign layer_0[125] = ~(in[132] ^ in[165]); 
    assign layer_0[126] = ~in[121] | (in[121] & in[163]); 
    assign layer_0[127] = in[164] & ~in[105]; 
    assign layer_0[128] = ~(in[117] | in[125]); 
    assign layer_0[129] = ~in[86] | (in[43] & in[86]); 
    assign layer_0[130] = in[37] | in[40]; 
    assign layer_0[131] = ~(in[36] | in[60]); 
    assign layer_0[132] = ~(in[232] | in[132]); 
    assign layer_0[133] = in[148] ^ in[235]; 
    assign layer_0[134] = ~in[28]; 
    assign layer_0[135] = ~in[182] | (in[182] & in[219]); 
    assign layer_0[136] = in[195] & ~in[45]; 
    assign layer_0[137] = in[227] ^ in[246]; 
    assign layer_0[138] = in[138] & ~in[171]; 
    assign layer_0[139] = ~(in[86] ^ in[22]); 
    assign layer_0[140] = in[135] ^ in[132]; 
    assign layer_0[141] = in[203] | in[108]; 
    assign layer_0[142] = in[164] | in[21]; 
    assign layer_0[143] = in[98] ^ in[102]; 
    assign layer_0[144] = ~(in[135] ^ in[228]); 
    assign layer_0[145] = in[82] ^ in[227]; 
    assign layer_0[146] = ~in[137]; 
    assign layer_0[147] = ~in[59] | (in[90] & in[59]); 
    assign layer_0[148] = ~(in[70] | in[54]); 
    assign layer_0[149] = ~(in[234] | in[28]); 
    assign layer_0[150] = in[163] | in[117]; 
    assign layer_0[151] = in[182] ^ in[229]; 
    assign layer_0[152] = ~in[24] | (in[24] & in[188]); 
    assign layer_0[153] = in[180] | in[212]; 
    assign layer_0[154] = in[214] | in[52]; 
    assign layer_0[155] = ~(in[119] | in[150]); 
    assign layer_0[156] = ~(in[201] ^ in[163]); 
    assign layer_0[157] = in[168] & ~in[162]; 
    assign layer_0[158] = ~(in[155] | in[171]); 
    assign layer_0[159] = in[39] | in[107]; 
    assign layer_0[160] = in[218] | in[103]; 
    assign layer_0[161] = ~(in[219] | in[44]); 
    assign layer_0[162] = ~(in[116] | in[114]); 
    assign layer_0[163] = in[124]; 
    assign layer_0[164] = in[154] ^ in[71]; 
    assign layer_0[165] = ~in[168] | (in[195] & in[168]); 
    assign layer_0[166] = ~(in[233] ^ in[58]); 
    assign layer_0[167] = in[214]; 
    assign layer_0[168] = in[111] | in[232]; 
    assign layer_0[169] = ~in[108]; 
    assign layer_0[170] = ~in[131] | (in[215] & in[131]); 
    assign layer_0[171] = in[171] & ~in[142]; 
    assign layer_0[172] = in[123] ^ in[61]; 
    assign layer_0[173] = ~in[108]; 
    assign layer_0[174] = ~(in[68] | in[181]); 
    assign layer_0[175] = in[115] | in[151]; 
    assign layer_0[176] = in[40] | in[181]; 
    assign layer_0[177] = ~(in[83] ^ in[52]); 
    assign layer_0[178] = in[230] ^ in[182]; 
    assign layer_0[179] = ~(in[78] | in[110]); 
    assign layer_0[180] = in[147]; 
    assign layer_0[181] = ~(in[249] | in[244]); 
    assign layer_0[182] = ~(in[183] ^ in[68]); 
    assign layer_0[183] = ~in[69] | (in[102] & in[69]); 
    assign layer_0[184] = ~(in[105] | in[105]); 
    assign layer_0[185] = in[102] & ~in[188]; 
    assign layer_0[186] = ~in[115]; 
    assign layer_0[187] = ~in[147] | (in[147] & in[210]); 
    assign layer_0[188] = in[123] | in[125]; 
    assign layer_0[189] = ~in[201] | (in[140] & in[201]); 
    assign layer_0[190] = in[170] | in[154]; 
    assign layer_0[191] = ~(in[133] | in[115]); 
    assign layer_0[192] = in[117] ^ in[85]; 
    assign layer_0[193] = in[109] | in[118]; 
    assign layer_0[194] = in[235] | in[149]; 
    assign layer_0[195] = ~(in[77] | in[51]); 
    assign layer_0[196] = ~in[197] | (in[227] & in[197]); 
    assign layer_0[197] = ~(in[91] | in[88]); 
    assign layer_0[198] = ~in[69] | (in[116] & in[69]); 
    assign layer_0[199] = in[92]; 
    assign layer_0[200] = ~(in[166] | in[102]); 
    assign layer_0[201] = ~(in[219] | in[233]); 
    assign layer_0[202] = ~(in[42] | in[135]); 
    assign layer_0[203] = ~(in[66] ^ in[217]); 
    assign layer_0[204] = in[179] ^ in[211]; 
    assign layer_0[205] = in[89] & ~in[108]; 
    assign layer_0[206] = in[108] ^ in[227]; 
    assign layer_0[207] = in[88] & ~in[84]; 
    assign layer_0[208] = ~(in[93] ^ in[75]); 
    assign layer_0[209] = in[25] ^ in[148]; 
    assign layer_0[210] = in[204] | in[203]; 
    assign layer_0[211] = in[150] & ~in[212]; 
    assign layer_0[212] = in[55] & in[138]; 
    assign layer_0[213] = ~(in[55] | in[60]); 
    assign layer_0[214] = in[185]; 
    assign layer_0[215] = in[179] ^ in[149]; 
    assign layer_0[216] = in[179] ^ in[213]; 
    assign layer_0[217] = ~(in[156] & in[186]); 
    assign layer_0[218] = ~(in[233] | in[52]); 
    assign layer_0[219] = ~in[121] | (in[25] & in[121]); 
    assign layer_0[220] = ~in[140]; 
    assign layer_0[221] = in[117] ^ in[103]; 
    assign layer_0[222] = ~in[216] | (in[216] & in[196]); 
    assign layer_0[223] = ~(in[186] | in[53]); 
    assign layer_0[224] = ~(in[68] ^ in[38]); 
    assign layer_0[225] = in[155]; 
    assign layer_0[226] = in[213] | in[94]; 
    assign layer_0[227] = in[247] | in[246]; 
    assign layer_0[228] = in[104] & ~in[101]; 
    assign layer_0[229] = in[231] ^ in[218]; 
    assign layer_0[230] = ~(in[26] | in[86]); 
    assign layer_0[231] = in[72] & in[122]; 
    assign layer_0[232] = ~(in[72] ^ in[67]); 
    assign layer_0[233] = in[87] ^ in[101]; 
    assign layer_0[234] = in[184] | in[162]; 
    assign layer_0[235] = ~(in[166] | in[164]); 
    assign layer_0[236] = in[53] ^ in[86]; 
    assign layer_0[237] = in[139] | in[124]; 
    assign layer_0[238] = ~(in[51] | in[84]); 
    assign layer_0[239] = ~(in[116] | in[169]); 
    assign layer_0[240] = in[202] ^ in[179]; 
    assign layer_0[241] = ~in[101] | (in[172] & in[101]); 
    assign layer_0[242] = in[141] ^ in[77]; 
    assign layer_0[243] = ~in[147] | (in[135] & in[147]); 
    assign layer_0[244] = ~in[201] | (in[201] & in[24]); 
    assign layer_0[245] = ~(in[139] | in[141]); 
    assign layer_0[246] = in[40] ^ in[196]; 
    assign layer_0[247] = ~(in[115] | in[219]); 
    assign layer_0[248] = ~(in[117] & in[101]); 
    assign layer_0[249] = ~in[104]; 
    assign layer_0[250] = in[229]; 
    assign layer_0[251] = in[217] ^ in[58]; 
    assign layer_0[252] = in[195]; 
    assign layer_0[253] = ~in[150] | (in[116] & in[150]); 
    assign layer_0[254] = in[109] ^ in[213]; 
    assign layer_0[255] = in[245] ^ in[214]; 
    assign layer_0[256] = in[82] | in[165]; 
    assign layer_0[257] = ~(in[234] | in[109]); 
    assign layer_0[258] = in[201] | in[130]; 
    assign layer_0[259] = in[83] ^ in[54]; 
    assign layer_0[260] = ~in[119] | (in[119] & in[101]); 
    assign layer_0[261] = in[42] & ~in[106]; 
    assign layer_0[262] = ~(in[67] ^ in[85]); 
    assign layer_0[263] = in[76] | in[59]; 
    assign layer_0[264] = in[167] | in[219]; 
    assign layer_0[265] = ~(in[180] | in[196]); 
    assign layer_0[266] = ~(in[58] ^ in[56]); 
    assign layer_0[267] = in[102] ^ in[99]; 
    assign layer_0[268] = ~(in[115] | in[45]); 
    assign layer_0[269] = in[78] | in[36]; 
    assign layer_0[270] = in[233] ^ in[124]; 
    assign layer_0[271] = ~(in[163] | in[182]); 
    assign layer_0[272] = in[167] | in[164]; 
    assign layer_0[273] = in[167]; 
    assign layer_0[274] = ~in[60] | (in[57] & in[60]); 
    assign layer_0[275] = in[162] | in[198]; 
    assign layer_0[276] = ~in[103] | (in[82] & in[103]); 
    assign layer_0[277] = ~(in[37] | in[138]); 
    assign layer_0[278] = ~(in[124] ^ in[158]); 
    assign layer_0[279] = in[124] | in[243]; 
    assign layer_0[280] = ~(in[155] | in[166]); 
    assign layer_0[281] = ~(in[180] ^ in[188]); 
    assign layer_0[282] = in[58]; 
    assign layer_0[283] = in[108] | in[54]; 
    assign layer_0[284] = in[131] ^ in[133]; 
    assign layer_0[285] = in[98] ^ in[186]; 
    assign layer_0[286] = in[172] | in[45]; 
    assign layer_0[287] = in[67] | in[123]; 
    assign layer_0[288] = in[186] & ~in[65]; 
    assign layer_0[289] = in[86] & ~in[204]; 
    assign layer_0[290] = in[185]; 
    assign layer_0[291] = in[244] | in[81]; 
    assign layer_0[292] = ~(in[36] ^ in[84]); 
    assign layer_0[293] = ~(in[148] ^ in[89]); 
    assign layer_0[294] = ~in[105] | (in[77] & in[105]); 
    assign layer_0[295] = in[168] | in[165]; 
    assign layer_0[296] = in[180] ^ in[89]; 
    assign layer_0[297] = ~(in[116] & in[156]); 
    assign layer_0[298] = ~(in[134] ^ in[25]); 
    assign layer_0[299] = ~in[57]; 
    assign layer_0[300] = in[163] ^ in[157]; 
    assign layer_0[301] = ~(in[180] ^ in[211]); 
    assign layer_0[302] = ~in[57] | (in[43] & in[57]); 
    assign layer_0[303] = ~(in[124] | in[42]); 
    assign layer_0[304] = in[130] ^ in[86]; 
    assign layer_0[305] = ~in[165]; 
    assign layer_0[306] = ~(in[140] & in[122]); 
    assign layer_0[307] = ~(in[105] ^ in[107]); 
    assign layer_0[308] = ~(in[187] | in[131]); 
    assign layer_0[309] = in[101] ^ in[99]; 
    assign layer_0[310] = in[198] & ~in[23]; 
    assign layer_0[311] = in[141] ^ in[188]; 
    assign layer_0[312] = ~(in[121] | in[116]); 
    assign layer_0[313] = ~(in[201] | in[185]); 
    assign layer_0[314] = in[198] & ~in[43]; 
    assign layer_0[315] = in[156] ^ in[202]; 
    assign layer_0[316] = ~in[170] | (in[170] & in[151]); 
    assign layer_0[317] = in[229] ^ in[51]; 
    assign layer_0[318] = in[165] ^ in[83]; 
    assign layer_0[319] = in[201] | in[217]; 
    assign layer_0[320] = in[178] | in[211]; 
    assign layer_0[321] = in[132] ^ in[150]; 
    assign layer_0[322] = ~in[132] | (in[132] & in[211]); 
    assign layer_0[323] = ~(in[110] | in[52]); 
    assign layer_0[324] = ~(in[169] ^ in[155]); 
    assign layer_0[325] = in[92] ^ in[123]; 
    assign layer_0[326] = in[226] ^ in[148]; 
    assign layer_0[327] = in[169] & ~in[197]; 
    assign layer_0[328] = ~(in[82] ^ in[104]); 
    assign layer_0[329] = ~(in[40] ^ in[87]); 
    assign layer_0[330] = ~(in[116] | in[86]); 
    assign layer_0[331] = in[167] ^ in[119]; 
    assign layer_0[332] = in[92]; 
    assign layer_0[333] = ~(in[142] | in[104]); 
    assign layer_0[334] = in[51]; 
    assign layer_0[335] = ~(in[92] | in[74]); 
    assign layer_0[336] = ~(in[132] ^ in[118]); 
    assign layer_0[337] = ~(in[89] ^ in[97]); 
    assign layer_0[338] = in[74] & ~in[156]; 
    assign layer_0[339] = in[195] | in[187]; 
    assign layer_0[340] = ~(in[116] ^ in[102]); 
    assign layer_0[341] = in[125] & ~in[137]; 
    assign layer_0[342] = ~(in[156] ^ in[203]); 
    assign layer_0[343] = ~in[201] | (in[108] & in[201]); 
    assign layer_0[344] = in[92] | in[212]; 
    assign layer_0[345] = ~(in[102] | in[220]); 
    assign layer_0[346] = ~(in[106] ^ in[134]); 
    assign layer_0[347] = in[85] ^ in[103]; 
    assign layer_0[348] = ~in[179]; 
    assign layer_0[349] = ~(in[201] ^ in[164]); 
    assign layer_0[350] = in[72] | in[83]; 
    assign layer_0[351] = in[220] | in[102]; 
    assign layer_0[352] = in[218] ^ in[185]; 
    assign layer_0[353] = ~in[105] | (in[82] & in[105]); 
    assign layer_0[354] = ~in[167] | (in[167] & in[226]); 
    assign layer_0[355] = in[184] & ~in[88]; 
    assign layer_0[356] = in[228] ^ in[166]; 
    assign layer_0[357] = ~in[135]; 
    assign layer_0[358] = ~(in[106] ^ in[75]); 
    assign layer_0[359] = ~(in[72] ^ in[54]); 
    assign layer_0[360] = in[61] ^ in[43]; 
    assign layer_0[361] = in[70] & ~in[62]; 
    assign layer_0[362] = in[104]; 
    assign layer_0[363] = in[93] | in[137]; 
    assign layer_0[364] = ~in[155]; 
    assign layer_0[365] = ~in[149] | (in[149] & in[229]); 
    assign layer_0[366] = ~(in[182] | in[131]); 
    assign layer_0[367] = in[40] | in[58]; 
    assign layer_0[368] = in[39] ^ in[22]; 
    assign layer_0[369] = in[216] & ~in[75]; 
    assign layer_0[370] = ~in[138]; 
    assign layer_0[371] = ~(in[57] ^ in[105]); 
    assign layer_0[372] = ~in[155] | (in[78] & in[155]); 
    assign layer_0[373] = ~(in[70] ^ in[86]); 
    assign layer_0[374] = in[152] ^ in[186]; 
    assign layer_0[375] = ~(in[246] ^ in[116]); 
    assign layer_0[376] = ~in[201] | (in[39] & in[201]); 
    assign layer_0[377] = in[135] & ~in[181]; 
    assign layer_0[378] = ~in[139]; 
    assign layer_0[379] = in[88] & ~in[59]; 
    assign layer_0[380] = ~(in[196] | in[217]); 
    assign layer_0[381] = ~(in[214] ^ in[203]); 
    assign layer_0[382] = in[133] ^ in[148]; 
    assign layer_0[383] = in[103] | in[94]; 
    assign layer_0[384] = ~(in[120] ^ in[95]); 
    assign layer_0[385] = ~(in[77] ^ in[56]); 
    assign layer_0[386] = ~(in[38] | in[187]); 
    assign layer_0[387] = in[187] & ~in[233]; 
    assign layer_0[388] = in[40] ^ in[54]; 
    assign layer_0[389] = ~in[164] | (in[229] & in[164]); 
    assign layer_0[390] = in[135] & in[134]; 
    assign layer_0[391] = in[135] & ~in[147]; 
    assign layer_0[392] = in[165] & ~in[147]; 
    assign layer_0[393] = in[100] ^ in[105]; 
    assign layer_0[394] = in[151] & in[150]; 
    assign layer_0[395] = in[87] ^ in[52]; 
    assign layer_0[396] = in[167] ^ in[149]; 
    assign layer_0[397] = in[57] | in[195]; 
    assign layer_0[398] = in[76] | in[154]; 
    assign layer_0[399] = in[168] ^ in[76]; 
    assign layer_0[400] = in[117] ^ in[114]; 
    assign layer_0[401] = in[216] & ~in[131]; 
    assign layer_0[402] = ~(in[156] ^ in[179]); 
    assign layer_0[403] = ~(in[218] ^ in[110]); 
    assign layer_0[404] = in[149] ^ in[141]; 
    assign layer_0[405] = ~(in[102] | in[132]); 
    assign layer_0[406] = ~(in[227] ^ in[151]); 
    assign layer_0[407] = in[122] & ~in[92]; 
    assign layer_0[408] = in[69] & in[134]; 
    assign layer_0[409] = ~(in[134] ^ in[113]); 
    assign layer_0[410] = in[180] & ~in[232]; 
    assign layer_0[411] = ~(in[90] ^ in[42]); 
    assign layer_0[412] = ~(in[57] ^ in[104]); 
    assign layer_0[413] = in[153]; 
    assign layer_0[414] = ~(in[117] ^ in[115]); 
    assign layer_0[415] = ~(in[127] | in[76]); 
    assign layer_0[416] = in[248] | in[251]; 
    assign layer_0[417] = ~in[184] | (in[184] & in[124]); 
    assign layer_0[418] = in[195] | in[186]; 
    assign layer_0[419] = in[25] | in[43]; 
    assign layer_0[420] = ~(in[204] | in[152]); 
    assign layer_0[421] = ~(in[228] | in[115]); 
    assign layer_0[422] = ~(in[178] | in[122]); 
    assign layer_0[423] = ~(in[196] ^ in[199]); 
    assign layer_0[424] = ~in[102] | (in[102] & in[23]); 
    assign layer_0[425] = in[169]; 
    assign layer_0[426] = ~(in[43] | in[135]); 
    assign layer_0[427] = ~in[70] | (in[37] & in[70]); 
    assign layer_0[428] = in[115] | in[226]; 
    assign layer_0[429] = in[101] ^ in[70]; 
    assign layer_0[430] = in[250] ^ in[46]; 
    assign layer_0[431] = ~(in[150] & in[215]); 
    assign layer_0[432] = ~(in[62] | in[55]); 
    assign layer_0[433] = in[114] | in[68]; 
    assign layer_0[434] = in[125] | in[67]; 
    assign layer_0[435] = ~in[168]; 
    assign layer_0[436] = in[71] & ~in[140]; 
    assign layer_0[437] = ~(in[231] ^ in[228]); 
    assign layer_0[438] = in[38] ^ in[198]; 
    assign layer_0[439] = in[82] | in[152]; 
    assign layer_0[440] = ~in[38] | (in[38] & in[84]); 
    assign layer_0[441] = in[69] | in[71]; 
    assign layer_0[442] = ~in[132]; 
    assign layer_0[443] = in[116] | in[91]; 
    assign layer_0[444] = ~(in[99] | in[58]); 
    assign layer_0[445] = in[42] ^ in[154]; 
    assign layer_0[446] = ~(in[181] ^ in[212]); 
    assign layer_0[447] = in[37] | in[173]; 
    assign layer_0[448] = in[85] ^ in[101]; 
    assign layer_0[449] = in[108] | in[109]; 
    assign layer_0[450] = ~(in[40] | in[76]); 
    assign layer_0[451] = ~in[69] | (in[69] & in[42]); 
    assign layer_0[452] = ~(in[164] | in[182]); 
    assign layer_0[453] = ~(in[165] | in[120]); 
    assign layer_0[454] = in[204] | in[116]; 
    assign layer_0[455] = ~in[153] | (in[179] & in[153]); 
    assign layer_0[456] = in[212] ^ in[86]; 
    assign layer_0[457] = in[85] & in[106]; 
    assign layer_0[458] = in[104] ^ in[85]; 
    assign layer_0[459] = ~(in[229] | in[246]); 
    assign layer_0[460] = ~(in[139] ^ in[134]); 
    assign layer_0[461] = in[119] & in[124]; 
    assign layer_0[462] = in[199] | in[141]; 
    assign layer_0[463] = ~in[200]; 
    assign layer_0[464] = in[154] ^ in[119]; 
    assign layer_0[465] = ~(in[159] | in[180]); 
    assign layer_0[466] = in[170] & ~in[124]; 
    assign layer_0[467] = in[139] ^ in[182]; 
    assign layer_0[468] = ~(in[101] | in[117]); 
    assign layer_0[469] = in[82] ^ in[140]; 
    assign layer_0[470] = in[42] | in[151]; 
    assign layer_0[471] = in[198] | in[178]; 
    assign layer_0[472] = ~(in[85] | in[115]); 
    assign layer_0[473] = in[131] ^ in[133]; 
    assign layer_0[474] = ~(in[148] & in[106]); 
    assign layer_0[475] = in[167] & ~in[234]; 
    assign layer_0[476] = ~(in[117] & in[133]); 
    assign layer_0[477] = ~(in[151] & in[182]); 
    assign layer_0[478] = ~in[174] | (in[174] & in[108]); 
    assign layer_0[479] = in[216] ^ in[167]; 
    assign layer_0[480] = ~(in[74] ^ in[99]); 
    assign layer_0[481] = ~in[229] | (in[229] & in[216]); 
    assign layer_0[482] = in[186] & in[57]; 
    assign layer_0[483] = ~in[120] | (in[120] & in[151]); 
    assign layer_0[484] = ~(in[105] ^ in[123]); 
    assign layer_0[485] = ~(in[147] | in[169]); 
    assign layer_0[486] = in[82] | in[51]; 
    assign layer_0[487] = ~(in[170] & in[167]); 
    assign layer_0[488] = ~(in[74] ^ in[107]); 
    assign layer_0[489] = ~(in[53] | in[26]); 
    assign layer_0[490] = ~(in[87] ^ in[69]); 
    assign layer_0[491] = ~in[165] | (in[84] & in[165]); 
    assign layer_0[492] = ~(in[104] ^ in[118]); 
    assign layer_0[493] = in[41] | in[73]; 
    assign layer_0[494] = in[117]; 
    assign layer_0[495] = in[140] | in[122]; 
    assign layer_0[496] = ~in[105]; 
    assign layer_0[497] = in[163] & ~in[85]; 
    assign layer_0[498] = in[182] | in[21]; 
    assign layer_0[499] = in[119] & in[120]; 
    assign layer_0[500] = ~(in[139] | in[108]); 
    assign layer_0[501] = in[166] & ~in[25]; 
    assign layer_0[502] = ~in[102] | (in[102] & in[39]); 
    assign layer_0[503] = ~(in[100] ^ in[69]); 
    assign layer_0[504] = ~(in[57] ^ in[109]); 
    assign layer_0[505] = ~(in[22] ^ in[114]); 
    assign layer_0[506] = in[186] ^ in[180]; 
    assign layer_0[507] = ~(in[124] | in[123]); 
    assign layer_0[508] = ~in[125] | (in[125] & in[136]); 
    assign layer_0[509] = ~(in[59] | in[37]); 
    assign layer_0[510] = in[251] | in[249]; 
    assign layer_0[511] = in[164] | in[249]; 
    assign layer_0[512] = ~(in[163] ^ in[105]); 
    assign layer_0[513] = in[197] & ~in[149]; 
    assign layer_0[514] = ~(in[78] | in[52]); 
    assign layer_0[515] = in[37] ^ in[102]; 
    assign layer_0[516] = in[216] | in[93]; 
    assign layer_0[517] = in[150] & in[165]; 
    assign layer_0[518] = in[105] & ~in[204]; 
    assign layer_0[519] = in[182] & ~in[99]; 
    assign layer_0[520] = ~(in[148] ^ in[166]); 
    assign layer_0[521] = ~in[89] | (in[76] & in[89]); 
    assign layer_0[522] = ~(in[229] | in[210]); 
    assign layer_0[523] = in[106] ^ in[138]; 
    assign layer_0[524] = ~(in[245] | in[127]); 
    assign layer_0[525] = in[135] & in[139]; 
    assign layer_0[526] = ~in[106]; 
    assign layer_0[527] = ~(in[122] ^ in[151]); 
    assign layer_0[528] = in[87] ^ in[84]; 
    assign layer_0[529] = ~(in[155] ^ in[121]); 
    assign layer_0[530] = in[115]; 
    assign layer_0[531] = in[51] | in[150]; 
    assign layer_0[532] = ~(in[36] | in[51]); 
    assign layer_0[533] = ~(in[124] | in[155]); 
    assign layer_0[534] = in[111] | in[215]; 
    assign layer_0[535] = in[105] & ~in[203]; 
    assign layer_0[536] = in[101] ^ in[115]; 
    assign layer_0[537] = ~(in[169] | in[110]); 
    assign layer_0[538] = ~(in[204] ^ in[124]); 
    assign layer_0[539] = ~(in[135] ^ in[165]); 
    assign layer_0[540] = ~(in[217] | in[186]); 
    assign layer_0[541] = in[109] | in[131]; 
    assign layer_0[542] = ~in[118] | (in[118] & in[173]); 
    assign layer_0[543] = ~(in[166] | in[131]); 
    assign layer_0[544] = ~(in[78] | in[105]); 
    assign layer_0[545] = in[150] | in[234]; 
    assign layer_0[546] = ~(in[61] ^ in[142]); 
    assign layer_0[547] = in[98] ^ in[140]; 
    assign layer_0[548] = ~(in[98] & in[102]); 
    assign layer_0[549] = in[42] ^ in[75]; 
    assign layer_0[550] = ~(in[107] | in[149]); 
    assign layer_0[551] = in[155]; 
    assign layer_0[552] = in[89]; 
    assign layer_0[553] = ~(in[139] | in[245]); 
    assign layer_0[554] = ~in[106]; 
    assign layer_0[555] = ~(in[24] | in[27]); 
    assign layer_0[556] = ~(in[142] ^ in[57]); 
    assign layer_0[557] = in[235] | in[140]; 
    assign layer_0[558] = ~(in[72] ^ in[43]); 
    assign layer_0[559] = in[125]; 
    assign layer_0[560] = ~(in[183] ^ in[163]); 
    assign layer_0[561] = ~in[86] | (in[86] & in[74]); 
    assign layer_0[562] = in[55] | in[86]; 
    assign layer_0[563] = in[133] ^ in[110]; 
    assign layer_0[564] = ~(in[181] ^ in[54]); 
    assign layer_0[565] = in[201] & ~in[154]; 
    assign layer_0[566] = ~in[37]; 
    assign layer_0[567] = ~(in[89] & in[90]); 
    assign layer_0[568] = in[84] ^ in[86]; 
    assign layer_0[569] = in[231] ^ in[120]; 
    assign layer_0[570] = ~(in[172] | in[139]); 
    assign layer_0[571] = ~(in[197] | in[24]); 
    assign layer_0[572] = in[199] & ~in[102]; 
    assign layer_0[573] = ~(in[233] ^ in[132]); 
    assign layer_0[574] = in[182] | in[164]; 
    assign layer_0[575] = ~(in[132] ^ in[27]); 
    assign layer_0[576] = in[227] ^ in[247]; 
    assign layer_0[577] = in[102] & ~in[73]; 
    assign layer_0[578] = ~in[60] | (in[148] & in[60]); 
    assign layer_0[579] = ~(in[167] ^ in[152]); 
    assign layer_0[580] = ~in[103] | (in[103] & in[92]); 
    assign layer_0[581] = in[132]; 
    assign layer_0[582] = in[124] | in[89]; 
    assign layer_0[583] = ~in[84] | (in[232] & in[84]); 
    assign layer_0[584] = ~(in[232] | in[200]); 
    assign layer_0[585] = in[188] | in[186]; 
    assign layer_0[586] = in[91] | in[204]; 
    assign layer_0[587] = in[26] | in[102]; 
    assign layer_0[588] = ~(in[110] | in[196]); 
    assign layer_0[589] = ~(in[117] | in[89]); 
    assign layer_0[590] = in[100] ^ in[102]; 
    assign layer_0[591] = ~in[184] | (in[87] & in[184]); 
    assign layer_0[592] = in[230] & ~in[181]; 
    assign layer_0[593] = in[181] | in[179]; 
    assign layer_0[594] = in[231] | in[215]; 
    assign layer_0[595] = ~in[133]; 
    assign layer_0[596] = ~(in[58] | in[75]); 
    assign layer_0[597] = ~(in[229] ^ in[197]); 
    assign layer_0[598] = in[40]; 
    assign layer_0[599] = in[87]; 
    assign layer_0[600] = ~in[53] | (in[53] & in[58]); 
    assign layer_0[601] = ~(in[102] | in[100]); 
    assign layer_0[602] = ~(in[54] ^ in[70]); 
    assign layer_0[603] = ~(in[26] | in[108]); 
    assign layer_0[604] = ~(in[170] | in[172]); 
    assign layer_0[605] = ~(in[123] | in[77]); 
    assign layer_0[606] = in[70] & ~in[201]; 
    assign layer_0[607] = in[109] | in[174]; 
    assign layer_0[608] = ~(in[237] ^ in[62]); 
    assign layer_0[609] = ~(in[197] ^ in[164]); 
    assign layer_0[610] = in[229] | in[68]; 
    assign layer_0[611] = in[42] ^ in[218]; 
    assign layer_0[612] = ~(in[140] ^ in[216]); 
    assign layer_0[613] = in[147] | in[107]; 
    assign layer_0[614] = in[106] ^ in[136]; 
    assign layer_0[615] = in[141] & in[173]; 
    assign layer_0[616] = ~(in[138] | in[44]); 
    assign layer_0[617] = ~(in[235] | in[169]); 
    assign layer_0[618] = in[169] ^ in[197]; 
    assign layer_0[619] = ~(in[141] | in[116]); 
    assign layer_0[620] = ~(in[91] ^ in[151]); 
    assign layer_0[621] = in[54] & ~in[100]; 
    assign layer_0[622] = in[248] | in[136]; 
    assign layer_0[623] = in[56] & ~in[228]; 
    assign layer_0[624] = in[135] & ~in[85]; 
    assign layer_0[625] = in[76] & ~in[73]; 
    assign layer_0[626] = ~(in[221] | in[99]); 
    assign layer_0[627] = in[140]; 
    assign layer_0[628] = ~in[150] | (in[233] & in[150]); 
    assign layer_0[629] = ~(in[154] | in[55]); 
    assign layer_0[630] = ~(in[77] | in[60]); 
    assign layer_0[631] = in[71] ^ in[212]; 
    assign layer_0[632] = in[105] & ~in[179]; 
    assign layer_0[633] = ~(in[246] ^ in[154]); 
    assign layer_0[634] = ~in[101] | (in[101] & in[24]); 
    assign layer_0[635] = in[77] | in[126]; 
    assign layer_0[636] = ~(in[131] | in[133]); 
    assign layer_0[637] = ~(in[147] | in[165]); 
    assign layer_0[638] = ~in[184] | (in[213] & in[184]); 
    assign layer_0[639] = in[198]; 
    assign layer_0[640] = ~(in[220] ^ in[189]); 
    assign layer_0[641] = ~in[106]; 
    assign layer_0[642] = in[214]; 
    assign layer_0[643] = in[199] & ~in[130]; 
    assign layer_0[644] = in[134] & ~in[125]; 
    assign layer_0[645] = ~(in[24] ^ in[117]); 
    assign layer_0[646] = ~(in[232] | in[67]); 
    assign layer_0[647] = in[120] | in[152]; 
    assign layer_0[648] = ~in[107] | (in[40] & in[107]); 
    assign layer_0[649] = in[122] ^ in[153]; 
    assign layer_0[650] = ~(in[153] ^ in[122]); 
    assign layer_0[651] = in[107] & ~in[155]; 
    assign layer_0[652] = in[69] | in[248]; 
    assign layer_0[653] = in[150] ^ in[123]; 
    assign layer_0[654] = ~(in[217] | in[218]); 
    assign layer_0[655] = ~(in[76] ^ in[70]); 
    assign layer_0[656] = in[58] | in[87]; 
    assign layer_0[657] = ~(in[108] ^ in[130]); 
    assign layer_0[658] = ~(in[138] ^ in[152]); 
    assign layer_0[659] = ~in[102] | (in[102] & in[211]); 
    assign layer_0[660] = in[133] & in[88]; 
    assign layer_0[661] = ~(in[109] | in[41]); 
    assign layer_0[662] = ~(in[88] ^ in[57]); 
    assign layer_0[663] = in[116] & ~in[231]; 
    assign layer_0[664] = ~(in[132] ^ in[150]); 
    assign layer_0[665] = ~in[86] | (in[74] & in[86]); 
    assign layer_0[666] = ~(in[92] ^ in[90]); 
    assign layer_0[667] = in[71]; 
    assign layer_0[668] = in[41] ^ in[74]; 
    assign layer_0[669] = ~(in[233] ^ in[150]); 
    assign layer_0[670] = ~(in[77] | in[167]); 
    assign layer_0[671] = ~in[75] | (in[75] & in[122]); 
    assign layer_0[672] = ~(in[76] ^ in[108]); 
    assign layer_0[673] = in[212] | in[214]; 
    assign layer_0[674] = in[52] ^ in[41]; 
    assign layer_0[675] = in[188] ^ in[178]; 
    assign layer_0[676] = ~(in[77] | in[108]); 
    assign layer_0[677] = ~(in[166] ^ in[147]); 
    assign layer_0[678] = in[73] & ~in[220]; 
    assign layer_0[679] = in[183] & ~in[90]; 
    assign layer_0[680] = in[196] ^ in[39]; 
    assign layer_0[681] = in[108] ^ in[140]; 
    assign layer_0[682] = ~in[104] | (in[172] & in[104]); 
    assign layer_0[683] = ~(in[24] ^ in[70]); 
    assign layer_0[684] = ~(in[170] ^ in[203]); 
    assign layer_0[685] = ~in[162] | (in[59] & in[162]); 
    assign layer_0[686] = ~in[39] | (in[39] & in[83]); 
    assign layer_0[687] = ~in[118] | (in[118] & in[199]); 
    assign layer_0[688] = ~in[51] | (in[51] & in[169]); 
    assign layer_0[689] = in[228] | in[85]; 
    assign layer_0[690] = in[150] & in[134]; 
    assign layer_0[691] = in[109] ^ in[42]; 
    assign layer_0[692] = in[86] & ~in[146]; 
    assign layer_0[693] = ~(in[150] ^ in[201]); 
    assign layer_0[694] = ~(in[70] ^ in[56]); 
    assign layer_0[695] = in[24] | in[156]; 
    assign layer_0[696] = in[149] ^ in[164]; 
    assign layer_0[697] = in[78] | in[142]; 
    assign layer_0[698] = in[150] | in[151]; 
    assign layer_0[699] = ~in[89] | (in[89] & in[54]); 
    assign layer_0[700] = ~(in[68] | in[99]); 
    assign layer_0[701] = ~(in[22] | in[94]); 
    assign layer_0[702] = in[154] | in[147]; 
    assign layer_0[703] = ~(in[150] | in[22]); 
    assign layer_0[704] = ~(in[229] ^ in[171]); 
    assign layer_0[705] = ~(in[116] | in[185]); 
    assign layer_0[706] = ~(in[41] | in[156]); 
    assign layer_0[707] = ~(in[231] | in[94]); 
    assign layer_0[708] = in[236] ^ in[250]; 
    assign layer_0[709] = ~(in[147] | in[205]); 
    assign layer_0[710] = in[182] & ~in[196]; 
    assign layer_0[711] = in[165] | in[102]; 
    assign layer_0[712] = in[153] ^ in[115]; 
    assign layer_0[713] = in[51] & in[220]; 
    assign layer_0[714] = ~in[166] | (in[166] & in[79]); 
    assign layer_0[715] = ~(in[109] | in[107]); 
    assign layer_0[716] = ~in[61]; 
    assign layer_0[717] = in[53] ^ in[83]; 
    assign layer_0[718] = ~(in[197] | in[189]); 
    assign layer_0[719] = ~(in[203] | in[216]); 
    assign layer_0[720] = in[71] | in[157]; 
    assign layer_0[721] = in[196] ^ in[227]; 
    assign layer_0[722] = ~(in[83] | in[91]); 
    assign layer_0[723] = ~in[43] | (in[43] & in[101]); 
    assign layer_0[724] = in[124] & ~in[216]; 
    assign layer_0[725] = ~(in[232] | in[115]); 
    assign layer_0[726] = ~(in[229] ^ in[21]); 
    assign layer_0[727] = in[38] ^ in[69]; 
    assign layer_0[728] = in[149] ^ in[55]; 
    assign layer_0[729] = ~(in[40] | in[37]); 
    assign layer_0[730] = in[180]; 
    assign layer_0[731] = ~(in[44] | in[40]); 
    assign layer_0[732] = in[135] | in[165]; 
    assign layer_0[733] = ~in[185] | (in[72] & in[185]); 
    assign layer_0[734] = in[198] ^ in[85]; 
    assign layer_0[735] = in[84] & ~in[92]; 
    assign layer_0[736] = in[230] ^ in[55]; 
    assign layer_0[737] = ~(in[78] | in[123]); 
    assign layer_0[738] = in[100] & ~in[41]; 
    assign layer_0[739] = ~in[123] | (in[42] & in[123]); 
    assign layer_0[740] = in[104] & ~in[60]; 
    assign layer_0[741] = in[203] | in[229]; 
    assign layer_0[742] = ~(in[57] | in[88]); 
    assign layer_0[743] = ~(in[84] ^ in[53]); 
    assign layer_0[744] = in[27] | in[54]; 
    assign layer_0[745] = in[150] ^ in[165]; 
    assign layer_0[746] = in[148] | in[166]; 
    assign layer_0[747] = in[151] & in[119]; 
    assign layer_0[748] = in[196] ^ in[228]; 
    assign layer_0[749] = in[72] & ~in[235]; 
    assign layer_0[750] = in[24] | in[195]; 
    assign layer_0[751] = in[197] | in[172]; 
    assign layer_0[752] = in[154] | in[246]; 
    assign layer_0[753] = in[87] ^ in[132]; 
    assign layer_0[754] = ~in[194] | (in[194] & in[156]); 
    assign layer_0[755] = in[150] ^ in[69]; 
    assign layer_0[756] = ~(in[132] ^ in[41]); 
    assign layer_0[757] = ~(in[149] ^ in[167]); 
    assign layer_0[758] = ~in[197] | (in[51] & in[197]); 
    assign layer_0[759] = ~(in[234] | in[166]); 
    assign layer_0[760] = ~(in[61] | in[99]); 
    assign layer_0[761] = in[117] & ~in[230]; 
    assign layer_0[762] = in[187] ^ in[181]; 
    assign layer_0[763] = in[170] | in[66]; 
    assign layer_0[764] = in[125] ^ in[149]; 
    assign layer_0[765] = in[104] & ~in[219]; 
    assign layer_0[766] = in[69] | in[116]; 
    assign layer_0[767] = ~(in[108] | in[189]); 
    assign layer_0[768] = in[92] & ~in[44]; 
    assign layer_0[769] = ~(in[100] ^ in[162]); 
    assign layer_0[770] = ~in[119] | (in[87] & in[119]); 
    assign layer_0[771] = in[51] | in[97]; 
    assign layer_0[772] = ~(in[156] | in[247]); 
    assign layer_0[773] = in[155] | in[44]; 
    assign layer_0[774] = ~(in[41] ^ in[43]); 
    assign layer_0[775] = ~(in[250] ^ in[57]); 
    assign layer_0[776] = ~(in[39] ^ in[53]); 
    assign layer_0[777] = ~(in[106] | in[109]); 
    assign layer_0[778] = ~in[88] | (in[181] & in[88]); 
    assign layer_0[779] = ~(in[217] | in[87]); 
    assign layer_0[780] = ~(in[184] | in[131]); 
    assign layer_0[781] = in[164] | in[166]; 
    assign layer_0[782] = ~in[119] | (in[113] & in[119]); 
    assign layer_0[783] = ~(in[72] ^ in[59]); 
    assign layer_0[784] = in[187] | in[141]; 
    assign layer_0[785] = ~in[73] | (in[203] & in[73]); 
    assign layer_0[786] = in[122]; 
    assign layer_0[787] = in[76]; 
    assign layer_0[788] = in[164] | in[187]; 
    assign layer_0[789] = in[44] | in[94]; 
    assign layer_0[790] = ~in[152] | (in[27] & in[152]); 
    assign layer_0[791] = ~in[148]; 
    assign layer_0[792] = ~(in[163] ^ in[170]); 
    assign layer_0[793] = in[234] ^ in[231]; 
    assign layer_0[794] = in[216] | in[188]; 
    assign layer_0[795] = ~(in[169] | in[200]); 
    assign layer_0[796] = ~(in[102] ^ in[219]); 
    assign layer_0[797] = in[84] ^ in[116]; 
    assign layer_0[798] = in[44] | in[221]; 
    assign layer_0[799] = in[188] | in[204]; 
    assign layer_0[800] = ~(in[204] ^ in[101]); 
    assign layer_0[801] = in[147] ^ in[165]; 
    assign layer_0[802] = ~(in[61] | in[94]); 
    assign layer_0[803] = ~(in[73] | in[83]); 
    assign layer_0[804] = ~(in[195] | in[168]); 
    assign layer_0[805] = ~(in[116] ^ in[134]); 
    assign layer_0[806] = in[132] | in[216]; 
    assign layer_0[807] = ~(in[106] ^ in[93]); 
    assign layer_0[808] = ~(in[198] ^ in[61]); 
    assign layer_0[809] = ~(in[60] | in[92]); 
    assign layer_0[810] = in[87] & ~in[178]; 
    assign layer_0[811] = in[73] | in[143]; 
    assign layer_0[812] = in[163] | in[118]; 
    assign layer_0[813] = in[227] | in[42]; 
    assign layer_0[814] = ~(in[205] ^ in[235]); 
    assign layer_0[815] = in[230] ^ in[217]; 
    assign layer_0[816] = in[186] ^ in[120]; 
    assign layer_0[817] = ~(in[119] | in[103]); 
    assign layer_0[818] = ~(in[202] | in[220]); 
    assign layer_0[819] = in[121] | in[137]; 
    assign layer_0[820] = ~in[147] | (in[135] & in[147]); 
    assign layer_0[821] = ~(in[150] & in[151]); 
    assign layer_0[822] = ~(in[186] & in[157]); 
    assign layer_0[823] = ~in[72] | (in[42] & in[72]); 
    assign layer_0[824] = ~(in[89] ^ in[92]); 
    assign layer_0[825] = in[124] ^ in[93]; 
    assign layer_0[826] = ~in[120] | (in[120] & in[188]); 
    assign layer_0[827] = in[99] ^ in[56]; 
    assign layer_0[828] = in[167] | in[66]; 
    assign layer_0[829] = ~(in[58] ^ in[89]); 
    assign layer_0[830] = ~(in[182] ^ in[196]); 
    assign layer_0[831] = ~in[94]; 
    assign layer_0[832] = ~in[100] | (in[100] & in[82]); 
    assign layer_0[833] = ~(in[71] | in[55]); 
    assign layer_0[834] = ~(in[178] | in[197]); 
    assign layer_0[835] = ~(in[166] ^ in[135]); 
    assign layer_0[836] = in[167]; 
    assign layer_0[837] = ~(in[216] | in[201]); 
    assign layer_0[838] = in[59] | in[55]; 
    assign layer_0[839] = in[36] | in[174]; 
    assign layer_0[840] = in[198] ^ in[228]; 
    assign layer_0[841] = ~in[70] | (in[37] & in[70]); 
    assign layer_0[842] = in[100] & ~in[88]; 
    assign layer_0[843] = in[198] | in[179]; 
    assign layer_0[844] = ~in[71] | (in[71] & in[136]); 
    assign layer_0[845] = ~(in[93] & in[123]); 
    assign layer_0[846] = in[62] ^ in[139]; 
    assign layer_0[847] = ~(in[54] ^ in[179]); 
    assign layer_0[848] = in[44] ^ in[77]; 
    assign layer_0[849] = in[55]; 
    assign layer_0[850] = ~in[110] | (in[139] & in[110]); 
    assign layer_0[851] = in[166]; 
    assign layer_0[852] = ~in[39] | (in[84] & in[39]); 
    assign layer_0[853] = ~in[216] | (in[216] & in[140]); 
    assign layer_0[854] = ~(in[183] ^ in[101]); 
    assign layer_0[855] = in[220] | in[111]; 
    assign layer_0[856] = ~(in[184] ^ in[52]); 
    assign layer_0[857] = ~(in[135] ^ in[247]); 
    assign layer_0[858] = in[217] | in[185]; 
    assign layer_0[859] = in[153] | in[23]; 
    assign layer_0[860] = ~(in[124] | in[107]); 
    assign layer_0[861] = ~in[198] | (in[198] & in[122]); 
    assign layer_0[862] = in[202] ^ in[155]; 
    assign layer_0[863] = ~(in[236] | in[116]); 
    assign layer_0[864] = in[24]; 
    assign layer_0[865] = ~(in[147] | in[203]); 
    assign layer_0[866] = ~(in[24] | in[195]); 
    assign layer_0[867] = in[164] ^ in[217]; 
    assign layer_0[868] = ~(in[107] ^ in[109]); 
    assign layer_0[869] = in[28]; 
    assign layer_0[870] = ~(in[228] ^ in[246]); 
    assign layer_0[871] = ~in[121] | (in[124] & in[121]); 
    assign layer_0[872] = ~in[148] | (in[150] & in[148]); 
    assign layer_0[873] = in[197] & ~in[151]; 
    assign layer_0[874] = ~(in[119] ^ in[93]); 
    assign layer_0[875] = in[166] ^ in[198]; 
    assign layer_0[876] = ~(in[228] | in[135]); 
    assign layer_0[877] = in[199] & ~in[26]; 
    assign layer_0[878] = ~in[119] | (in[119] & in[172]); 
    assign layer_0[879] = ~(in[99] ^ in[68]); 
    assign layer_0[880] = in[24] ^ in[170]; 
    assign layer_0[881] = in[101] | in[109]; 
    assign layer_0[882] = ~in[119] | (in[99] & in[119]); 
    assign layer_0[883] = ~(in[21] ^ in[23]); 
    assign layer_0[884] = in[169] ^ in[44]; 
    assign layer_0[885] = ~(in[181] ^ in[149]); 
    assign layer_0[886] = ~(in[90] | in[92]); 
    assign layer_0[887] = ~(in[197] ^ in[93]); 
    assign layer_0[888] = ~in[90] | (in[135] & in[90]); 
    assign layer_0[889] = in[204] ^ in[62]; 
    assign layer_0[890] = in[147] ^ in[181]; 
    assign layer_0[891] = in[213] ^ in[150]; 
    assign layer_0[892] = in[118] ^ in[130]; 
    assign layer_0[893] = ~in[104] | (in[104] & in[76]); 
    assign layer_0[894] = in[75] ^ in[131]; 
    assign layer_0[895] = in[166] & ~in[157]; 
    assign layer_0[896] = in[182] & ~in[58]; 
    assign layer_0[897] = in[126] & ~in[108]; 
    assign layer_0[898] = ~(in[124] | in[59]); 
    assign layer_0[899] = ~(in[23] | in[180]); 
    assign layer_0[900] = ~(in[190] | in[116]); 
    assign layer_0[901] = in[150] & ~in[126]; 
    assign layer_0[902] = ~in[199] | (in[164] & in[199]); 
    assign layer_0[903] = in[29] | in[87]; 
    assign layer_0[904] = in[152] ^ in[212]; 
    assign layer_0[905] = ~(in[185] ^ in[124]); 
    assign layer_0[906] = ~in[148]; 
    assign layer_0[907] = in[44]; 
    assign layer_0[908] = in[148] | in[56]; 
    assign layer_0[909] = ~(in[41] ^ in[106]); 
    assign layer_0[910] = ~(in[116] | in[57]); 
    assign layer_0[911] = ~(in[43] ^ in[25]); 
    assign layer_0[912] = ~(in[88] ^ in[212]); 
    assign layer_0[913] = in[77] | in[109]; 
    assign layer_0[914] = ~(in[141] & in[131]); 
    assign layer_0[915] = in[134] & ~in[204]; 
    assign layer_0[916] = ~(in[147] ^ in[133]); 
    assign layer_0[917] = ~(in[197] & in[118]); 
    assign layer_0[918] = in[148] & ~in[37]; 
    assign layer_0[919] = ~(in[167] ^ in[120]); 
    assign layer_0[920] = ~(in[217] & in[167]); 
    assign layer_0[921] = ~(in[188] ^ in[215]); 
    assign layer_0[922] = in[234] | in[201]; 
    assign layer_0[923] = in[248] ^ in[125]; 
    assign layer_0[924] = in[25] ^ in[85]; 
    assign layer_0[925] = ~in[199] | (in[37] & in[199]); 
    assign layer_0[926] = in[24] ^ in[226]; 
    assign layer_0[927] = in[155] ^ in[186]; 
    assign layer_0[928] = in[73] ^ in[103]; 
    assign layer_0[929] = ~(in[83] | in[148]); 
    assign layer_0[930] = in[202] ^ in[171]; 
    assign layer_0[931] = in[136]; 
    assign layer_0[932] = in[197] & ~in[84]; 
    assign layer_0[933] = ~(in[118] ^ in[132]); 
    assign layer_0[934] = ~(in[154] ^ in[123]); 
    assign layer_0[935] = in[219]; 
    assign layer_0[936] = ~(in[149] | in[147]); 
    assign layer_0[937] = ~(in[180] ^ in[183]); 
    assign layer_0[938] = in[196] | in[150]; 
    assign layer_0[939] = in[152] | in[82]; 
    assign layer_0[940] = ~(in[72] & in[121]); 
    assign layer_0[941] = in[102] | in[201]; 
    assign layer_0[942] = in[140] ^ in[91]; 
    assign layer_0[943] = ~(in[56] | in[92]); 
    assign layer_0[944] = ~(in[170] | in[171]); 
    assign layer_0[945] = in[40] ^ in[170]; 
    assign layer_0[946] = ~(in[54] | in[107]); 
    assign layer_0[947] = ~(in[148] | in[165]); 
    assign layer_0[948] = in[123] & ~in[212]; 
    assign layer_0[949] = in[125] | in[108]; 
    assign layer_0[950] = in[200] ^ in[233]; 
    assign layer_0[951] = ~(in[218] | in[123]); 
    assign layer_0[952] = in[218] | in[86]; 
    assign layer_0[953] = ~(in[180] ^ in[216]); 
    assign layer_0[954] = ~(in[82] | in[73]); 
    assign layer_0[955] = ~in[153]; 
    assign layer_0[956] = ~(in[186] | in[155]); 
    assign layer_0[957] = in[234] | in[220]; 
    assign layer_0[958] = in[162] ^ in[185]; 
    assign layer_0[959] = ~(in[148] ^ in[200]); 
    assign layer_0[960] = ~in[88]; 
    assign layer_0[961] = ~(in[120] ^ in[166]); 
    assign layer_0[962] = ~(in[210] | in[230]); 
    assign layer_0[963] = ~(in[183] ^ in[197]); 
    assign layer_0[964] = ~in[107] | (in[107] & in[157]); 
    assign layer_0[965] = in[120]; 
    assign layer_0[966] = ~(in[219] | in[136]); 
    assign layer_0[967] = ~(in[124] | in[149]); 
    assign layer_0[968] = in[213] & in[215]; 
    assign layer_0[969] = ~(in[99] ^ in[117]); 
    assign layer_0[970] = in[139] ^ in[153]; 
    assign layer_0[971] = ~(in[228] ^ in[52]); 
    assign layer_0[972] = ~(in[232] ^ in[235]); 
    assign layer_0[973] = in[147]; 
    assign layer_0[974] = ~(in[149] | in[131]); 
    assign layer_0[975] = in[131] | in[53]; 
    assign layer_0[976] = in[147] | in[185]; 
    assign layer_0[977] = in[51] | in[179]; 
    assign layer_0[978] = in[134] & in[131]; 
    assign layer_0[979] = in[42] ^ in[142]; 
    assign layer_0[980] = in[148] | in[163]; 
    assign layer_0[981] = in[206]; 
    assign layer_0[982] = in[92] | in[71]; 
    assign layer_0[983] = ~(in[132] ^ in[134]); 
    assign layer_0[984] = ~in[132] | (in[132] & in[73]); 
    assign layer_0[985] = in[185] ^ in[71]; 
    assign layer_0[986] = in[108] ^ in[77]; 
    assign layer_0[987] = in[163] ^ in[149]; 
    assign layer_0[988] = ~in[119] | (in[50] & in[119]); 
    assign layer_0[989] = in[168] | in[107]; 
    assign layer_0[990] = in[87] ^ in[41]; 
    assign layer_0[991] = ~(in[181] ^ in[233]); 
    assign layer_0[992] = in[67] | in[213]; 
    assign layer_0[993] = ~in[73] | (in[173] & in[73]); 
    assign layer_0[994] = in[107] | in[69]; 
    assign layer_0[995] = in[116] ^ in[114]; 
    assign layer_0[996] = in[148] | in[119]; 
    assign layer_0[997] = in[69] & in[101]; 
    assign layer_0[998] = in[67]; 
    assign layer_0[999] = in[108]; 
    assign layer_0[1000] = in[158] ^ in[205]; 
    assign layer_0[1001] = in[198] | in[213]; 
    assign layer_0[1002] = ~(in[130] ^ in[230]); 
    assign layer_0[1003] = in[132] & ~in[111]; 
    assign layer_0[1004] = ~in[117] | (in[143] & in[117]); 
    assign layer_0[1005] = in[148] | in[162]; 
    assign layer_0[1006] = in[185] | in[203]; 
    assign layer_0[1007] = in[183]; 
    assign layer_0[1008] = in[114] | in[235]; 
    assign layer_0[1009] = ~(in[169] ^ in[84]); 
    assign layer_0[1010] = ~(in[42] | in[200]); 
    assign layer_0[1011] = in[218] | in[102]; 
    assign layer_0[1012] = in[139] & ~in[41]; 
    assign layer_0[1013] = ~in[146]; 
    assign layer_0[1014] = ~(in[172] ^ in[203]); 
    assign layer_0[1015] = ~(in[101] ^ in[67]); 
    assign layer_0[1016] = ~(in[84] | in[165]); 
    assign layer_0[1017] = ~in[120] | (in[120] & in[213]); 
    assign layer_0[1018] = in[121] ^ in[123]; 
    assign layer_0[1019] = ~(in[135] ^ in[150]); 
    assign layer_0[1020] = in[115]; 
    assign layer_0[1021] = ~(in[181] ^ in[212]); 
    assign layer_0[1022] = ~in[166]; 
    assign layer_0[1023] = in[150]; 
    assign layer_0[1024] = in[100] ^ in[133]; 
    assign layer_0[1025] = in[132] | in[131]; 
    assign layer_0[1026] = ~(in[226] | in[97]); 
    assign layer_0[1027] = in[171] ^ in[217]; 
    assign layer_0[1028] = ~in[133] | (in[250] & in[133]); 
    assign layer_0[1029] = ~(in[99] | in[86]); 
    assign layer_0[1030] = in[90] & ~in[92]; 
    assign layer_0[1031] = ~(in[233] ^ in[230]); 
    assign layer_0[1032] = ~in[204] | (in[231] & in[204]); 
    assign layer_0[1033] = in[171] ^ in[180]; 
    assign layer_0[1034] = in[90] ^ in[108]; 
    assign layer_0[1035] = ~(in[84] | in[57]); 
    assign layer_0[1036] = ~in[247]; 
    assign layer_0[1037] = in[170] & ~in[141]; 
    assign layer_0[1038] = in[156] ^ in[154]; 
    assign layer_0[1039] = ~(in[245] | in[154]); 
    assign layer_0[1040] = in[157] | in[43]; 
    assign layer_0[1041] = ~(in[52] | in[178]); 
    assign layer_0[1042] = in[197]; 
    assign layer_0[1043] = ~(in[94] | in[103]); 
    assign layer_0[1044] = in[108] | in[139]; 
    assign layer_0[1045] = in[55] & ~in[38]; 
    assign layer_0[1046] = ~in[88] | (in[198] & in[88]); 
    assign layer_0[1047] = ~(in[125] | in[219]); 
    assign layer_0[1048] = ~in[72] | (in[77] & in[72]); 
    assign layer_0[1049] = in[148] ^ in[204]; 
    assign layer_0[1050] = in[55] & ~in[57]; 
    assign layer_0[1051] = in[108]; 
    assign layer_0[1052] = ~in[137] | (in[137] & in[196]); 
    assign layer_0[1053] = in[40] ^ in[107]; 
    assign layer_0[1054] = ~in[231] | (in[231] & in[164]); 
    assign layer_0[1055] = in[142] ^ in[155]; 
    assign layer_0[1056] = ~(in[90] ^ in[93]); 
    assign layer_0[1057] = ~in[73] | (in[62] & in[73]); 
    assign layer_0[1058] = ~(in[230] ^ in[227]); 
    assign layer_0[1059] = in[154] ^ in[118]; 
    assign layer_0[1060] = in[103]; 
    assign layer_0[1061] = ~in[103] | (in[103] & in[83]); 
    assign layer_0[1062] = in[136] | in[182]; 
    assign layer_0[1063] = in[55] | in[178]; 
    assign layer_0[1064] = in[56] & ~in[227]; 
    assign layer_0[1065] = ~(in[196] ^ in[182]); 
    assign layer_0[1066] = in[61] | in[235]; 
    assign layer_0[1067] = in[57] & ~in[44]; 
    assign layer_0[1068] = in[101] ^ in[118]; 
    assign layer_0[1069] = in[72] | in[88]; 
    assign layer_0[1070] = in[100] ^ in[102]; 
    assign layer_0[1071] = in[67]; 
    assign layer_0[1072] = in[132] | in[227]; 
    assign layer_0[1073] = ~(in[162] | in[70]); 
    assign layer_0[1074] = ~(in[231] ^ in[228]); 
    assign layer_0[1075] = in[68] ^ in[134]; 
    assign layer_0[1076] = in[151] | in[154]; 
    assign layer_0[1077] = in[67] | in[249]; 
    assign layer_0[1078] = in[133] & ~in[158]; 
    assign layer_0[1079] = ~(in[179] ^ in[54]); 
    assign layer_0[1080] = in[90] & ~in[134]; 
    assign layer_0[1081] = ~(in[246] ^ in[228]); 
    assign layer_0[1082] = ~(in[213] | in[135]); 
    assign layer_0[1083] = in[166] & ~in[134]; 
    assign layer_0[1084] = ~(in[60] ^ in[92]); 
    assign layer_0[1085] = ~(in[231] | in[22]); 
    assign layer_0[1086] = ~in[70] | (in[70] & in[59]); 
    assign layer_0[1087] = ~(in[98] ^ in[72]); 
    assign layer_0[1088] = in[106] | in[76]; 
    assign layer_0[1089] = ~(in[92] | in[91]); 
    assign layer_0[1090] = in[122] | in[139]; 
    assign layer_0[1091] = ~(in[43] | in[233]); 
    assign layer_0[1092] = ~(in[109] | in[91]); 
    assign layer_0[1093] = in[43] ^ in[91]; 
    assign layer_0[1094] = ~in[90] | (in[90] & in[46]); 
    assign layer_0[1095] = in[111] | in[63]; 
    assign layer_0[1096] = in[149] & ~in[154]; 
    assign layer_0[1097] = ~(in[188] ^ in[185]); 
    assign layer_0[1098] = in[170] | in[139]; 
    assign layer_0[1099] = in[123] & ~in[170]; 
    assign layer_0[1100] = ~in[152]; 
    assign layer_0[1101] = ~(in[157] | in[155]); 
    assign layer_0[1102] = ~(in[202] | in[219]); 
    assign layer_0[1103] = ~(in[107] ^ in[39]); 
    assign layer_0[1104] = in[152] | in[108]; 
    assign layer_0[1105] = ~in[122] | (in[122] & in[220]); 
    assign layer_0[1106] = in[154] & ~in[52]; 
    assign layer_0[1107] = ~(in[43] | in[57]); 
    assign layer_0[1108] = in[89] ^ in[76]; 
    assign layer_0[1109] = in[118] ^ in[169]; 
    assign layer_0[1110] = ~(in[131] | in[149]); 
    assign layer_0[1111] = in[114] | in[74]; 
    assign layer_0[1112] = ~(in[133] ^ in[102]); 
    assign layer_0[1113] = ~(in[218] ^ in[187]); 
    assign layer_0[1114] = in[46] | in[124]; 
    assign layer_0[1115] = in[56] & ~in[172]; 
    assign layer_0[1116] = in[42] ^ in[171]; 
    assign layer_0[1117] = ~in[60]; 
    assign layer_0[1118] = in[154] ^ in[38]; 
    assign layer_0[1119] = in[154] & ~in[22]; 
    assign layer_0[1120] = ~(in[247] ^ in[91]); 
    assign layer_0[1121] = ~(in[92] ^ in[250]); 
    assign layer_0[1122] = ~(in[187] | in[102]); 
    assign layer_0[1123] = in[88] & ~in[71]; 
    assign layer_0[1124] = ~(in[120] & in[88]); 
    assign layer_0[1125] = in[85] | in[99]; 
    assign layer_0[1126] = ~(in[202] ^ in[181]); 
    assign layer_0[1127] = ~in[180] | (in[180] & in[203]); 
    assign layer_0[1128] = in[249] ^ in[137]; 
    assign layer_0[1129] = ~in[87] | (in[87] & in[121]); 
    assign layer_0[1130] = in[138]; 
    assign layer_0[1131] = in[125]; 
    assign layer_0[1132] = ~(in[107] | in[91]); 
    assign layer_0[1133] = ~in[186] | (in[186] & in[248]); 
    assign layer_0[1134] = ~in[153]; 
    assign layer_0[1135] = in[149] ^ in[69]; 
    assign layer_0[1136] = ~(in[94] ^ in[26]); 
    assign layer_0[1137] = ~in[121] | (in[155] & in[121]); 
    assign layer_0[1138] = in[109] ^ in[123]; 
    assign layer_0[1139] = ~(in[75] & in[185]); 
    assign layer_0[1140] = ~(in[154] | in[138]); 
    assign layer_0[1141] = ~(in[27] | in[45]); 
    assign layer_0[1142] = ~(in[204] | in[62]); 
    assign layer_0[1143] = in[92] | in[70]; 
    assign layer_0[1144] = ~in[57] | (in[57] & in[120]); 
    assign layer_0[1145] = ~in[217] | (in[214] & in[217]); 
    assign layer_0[1146] = ~(in[117] ^ in[134]); 
    assign layer_0[1147] = in[166] & ~in[110]; 
    assign layer_0[1148] = ~(in[89] ^ in[45]); 
    assign layer_0[1149] = in[83] | in[92]; 
    assign layer_0[1150] = in[122] & ~in[197]; 
    assign layer_0[1151] = in[250] | in[91]; 
    assign layer_0[1152] = ~(in[100] ^ in[117]); 
    assign layer_0[1153] = in[56]; 
    assign layer_0[1154] = in[85] | in[70]; 
    assign layer_0[1155] = in[146]; 
    assign layer_0[1156] = ~(in[85] ^ in[71]); 
    assign layer_0[1157] = ~(in[70] ^ in[73]); 
    assign layer_0[1158] = in[248] ^ in[215]; 
    assign layer_0[1159] = in[173] ^ in[203]; 
    assign layer_0[1160] = ~in[109] | (in[109] & in[127]); 
    assign layer_0[1161] = in[122] & ~in[90]; 
    assign layer_0[1162] = in[137] & ~in[146]; 
    assign layer_0[1163] = in[106]; 
    assign layer_0[1164] = ~(in[139] | in[61]); 
    assign layer_0[1165] = ~(in[117] ^ in[228]); 
    assign layer_0[1166] = ~(in[182] ^ in[229]); 
    assign layer_0[1167] = in[61] | in[217]; 
    assign layer_0[1168] = in[236] ^ in[108]; 
    assign layer_0[1169] = ~(in[56] ^ in[131]); 
    assign layer_0[1170] = in[183] ^ in[84]; 
    assign layer_0[1171] = ~in[117] | (in[117] & in[103]); 
    assign layer_0[1172] = ~(in[202] ^ in[195]); 
    assign layer_0[1173] = ~in[55]; 
    assign layer_0[1174] = in[109] | in[108]; 
    assign layer_0[1175] = in[230] ^ in[134]; 
    assign layer_0[1176] = ~(in[157] | in[155]); 
    assign layer_0[1177] = in[139] ^ in[170]; 
    assign layer_0[1178] = in[137] & in[151]; 
    assign layer_0[1179] = in[75] & ~in[83]; 
    assign layer_0[1180] = ~(in[189] ^ in[213]); 
    assign layer_0[1181] = ~(in[236] ^ in[228]); 
    assign layer_0[1182] = in[75] ^ in[99]; 
    assign layer_0[1183] = ~(in[60] ^ in[54]); 
    assign layer_0[1184] = ~(in[60] | in[75]); 
    assign layer_0[1185] = in[134] & ~in[180]; 
    assign layer_0[1186] = ~in[165] | (in[165] & in[195]); 
    assign layer_0[1187] = ~(in[133] & in[102]); 
    assign layer_0[1188] = ~(in[170] ^ in[67]); 
    assign layer_0[1189] = in[164] & in[213]; 
    assign layer_0[1190] = in[89] ^ in[52]; 
    assign layer_0[1191] = in[90] ^ in[53]; 
    assign layer_0[1192] = ~(in[250] ^ in[153]); 
    assign layer_0[1193] = ~(in[201] | in[162]); 
    assign layer_0[1194] = ~(in[156] ^ in[124]); 
    assign layer_0[1195] = in[201]; 
    assign layer_0[1196] = in[101] & ~in[166]; 
    assign layer_0[1197] = ~(in[38] | in[163]); 
    assign layer_0[1198] = in[174] ^ in[38]; 
    assign layer_0[1199] = in[166] & ~in[141]; 
    assign layer_0[1200] = ~in[108] | (in[122] & in[108]); 
    assign layer_0[1201] = in[75] ^ in[57]; 
    assign layer_0[1202] = ~(in[149] | in[147]); 
    assign layer_0[1203] = ~(in[201] ^ in[195]); 
    assign layer_0[1204] = in[36] | in[106]; 
    assign layer_0[1205] = ~in[91]; 
    assign layer_0[1206] = ~in[58]; 
    assign layer_0[1207] = ~(in[102] | in[100]); 
    assign layer_0[1208] = in[121] & ~in[219]; 
    assign layer_0[1209] = ~in[133]; 
    assign layer_0[1210] = ~in[183] | (in[183] & in[127]); 
    assign layer_0[1211] = in[154] | in[62]; 
    assign layer_0[1212] = ~(in[232] | in[247]); 
    assign layer_0[1213] = ~(in[148] | in[99]); 
    assign layer_0[1214] = in[171] & ~in[196]; 
    assign layer_0[1215] = in[211] ^ in[88]; 
    assign layer_0[1216] = in[116] ^ in[211]; 
    assign layer_0[1217] = in[115] ^ in[148]; 
    assign layer_0[1218] = ~(in[151] ^ in[149]); 
    assign layer_0[1219] = ~(in[163] ^ in[249]); 
    assign layer_0[1220] = ~(in[178] | in[230]); 
    assign layer_0[1221] = in[90] & ~in[78]; 
    assign layer_0[1222] = in[115]; 
    assign layer_0[1223] = in[165] ^ in[25]; 
    assign layer_0[1224] = in[133] & ~in[25]; 
    assign layer_0[1225] = in[40] & ~in[70]; 
    assign layer_0[1226] = ~(in[135] ^ in[148]); 
    assign layer_0[1227] = ~in[100] | (in[100] & in[134]); 
    assign layer_0[1228] = in[196] & ~in[98]; 
    assign layer_0[1229] = ~(in[161] | in[211]); 
    assign layer_0[1230] = ~in[151] | (in[141] & in[151]); 
    assign layer_0[1231] = ~(in[86] ^ in[39]); 
    assign layer_0[1232] = in[115] ^ in[133]; 
    assign layer_0[1233] = in[93] | in[122]; 
    assign layer_0[1234] = in[133] & in[134]; 
    assign layer_0[1235] = ~(in[83] | in[243]); 
    assign layer_0[1236] = in[197] | in[99]; 
    assign layer_0[1237] = ~in[170] | (in[122] & in[170]); 
    assign layer_0[1238] = in[182] ^ in[61]; 
    assign layer_0[1239] = ~(in[182] ^ in[188]); 
    assign layer_0[1240] = ~(in[45] ^ in[74]); 
    assign layer_0[1241] = in[74] | in[61]; 
    assign layer_0[1242] = in[123] ^ in[154]; 
    assign layer_0[1243] = in[77] & ~in[123]; 
    assign layer_0[1244] = in[138] ^ in[171]; 
    assign layer_0[1245] = in[137] | in[210]; 
    assign layer_0[1246] = in[43] ^ in[89]; 
    assign layer_0[1247] = in[91] ^ in[89]; 
    assign layer_0[1248] = in[119] | in[203]; 
    assign layer_0[1249] = in[216] ^ in[200]; 
    assign layer_0[1250] = ~(in[100] | in[98]); 
    assign layer_0[1251] = in[119]; 
    assign layer_0[1252] = in[164] ^ in[167]; 
    assign layer_0[1253] = in[103]; 
    assign layer_0[1254] = in[201] & ~in[53]; 
    assign layer_0[1255] = ~(in[168] & in[105]); 
    assign layer_0[1256] = in[99] ^ in[102]; 
    assign layer_0[1257] = in[197] ^ in[187]; 
    assign layer_0[1258] = ~(in[57] ^ in[58]); 
    assign layer_0[1259] = in[131] | in[101]; 
    assign layer_0[1260] = ~in[93] | (in[93] & in[210]); 
    assign layer_0[1261] = in[75] | in[218]; 
    assign layer_0[1262] = in[181] & ~in[130]; 
    assign layer_0[1263] = ~(in[86] | in[100]); 
    assign layer_0[1264] = in[196] | in[61]; 
    assign layer_0[1265] = in[58] & ~in[248]; 
    assign layer_0[1266] = in[167] & ~in[229]; 
    assign layer_0[1267] = in[179] | in[69]; 
    assign layer_0[1268] = in[155] & ~in[121]; 
    assign layer_0[1269] = in[56] ^ in[93]; 
    assign layer_0[1270] = in[99] | in[243]; 
    assign layer_0[1271] = ~(in[127] | in[195]); 
    assign layer_0[1272] = ~in[86] | (in[135] & in[86]); 
    assign layer_0[1273] = in[58] | in[74]; 
    assign layer_0[1274] = ~(in[115] | in[102]); 
    assign layer_0[1275] = ~in[60]; 
    assign layer_0[1276] = in[86] | in[93]; 
    assign layer_0[1277] = in[100] | in[98]; 
    assign layer_0[1278] = ~(in[74] | in[158]); 
    assign layer_0[1279] = in[197]; 
    // Layer 1 ============================================================
    assign out[0] = layer_0[149]; 
    assign out[1] = layer_0[289] & layer_0[462]; 
    assign out[2] = layer_0[1138]; 
    assign out[3] = layer_0[218] & ~layer_0[1245]; 
    assign out[4] = layer_0[710] | layer_0[1189]; 
    assign out[5] = layer_0[4] & ~layer_0[278]; 
    assign out[6] = layer_0[3] & ~layer_0[1202]; 
    assign out[7] = ~layer_0[507]; 
    assign out[8] = ~layer_0[122] | (layer_0[613] & layer_0[122]); 
    assign out[9] = ~(layer_0[678] ^ layer_0[1116]); 
    assign out[10] = ~layer_0[957]; 
    assign out[11] = ~(layer_0[651] | layer_0[411]); 
    assign out[12] = ~layer_0[159] | (layer_0[9] & layer_0[159]); 
    assign out[13] = layer_0[27] & layer_0[400]; 
    assign out[14] = ~layer_0[622]; 
    assign out[15] = layer_0[18] & ~layer_0[1059]; 
    assign out[16] = ~layer_0[480]; 
    assign out[17] = layer_0[1143] & ~layer_0[844]; 
    assign out[18] = layer_0[211]; 
    assign out[19] = layer_0[642] ^ layer_0[0]; 
    assign out[20] = layer_0[877] & ~layer_0[803]; 
    assign out[21] = layer_0[225] & layer_0[761]; 
    assign out[22] = layer_0[144] & ~layer_0[322]; 
    assign out[23] = ~(layer_0[328] ^ layer_0[955]); 
    assign out[24] = ~(layer_0[705] | layer_0[974]); 
    assign out[25] = layer_0[843]; 
    assign out[26] = layer_0[49]; 
    assign out[27] = ~layer_0[989] | (layer_0[989] & layer_0[514]); 
    assign out[28] = ~(layer_0[872] | layer_0[741]); 
    assign out[29] = ~(layer_0[498] ^ layer_0[1221]); 
    assign out[30] = layer_0[973] & layer_0[607]; 
    assign out[31] = layer_0[1145] & ~layer_0[305]; 
    assign out[32] = layer_0[919]; 
    assign out[33] = layer_0[76] & ~layer_0[1278]; 
    assign out[34] = layer_0[806]; 
    assign out[35] = ~(layer_0[372] ^ layer_0[793]); 
    assign out[36] = layer_0[976]; 
    assign out[37] = ~(layer_0[872] | layer_0[393]); 
    assign out[38] = ~(layer_0[1233] ^ layer_0[1030]); 
    assign out[39] = layer_0[516]; 
    assign out[40] = ~layer_0[377]; 
    assign out[41] = layer_0[219] & ~layer_0[1107]; 
    assign out[42] = ~(layer_0[661] & layer_0[190]); 
    assign out[43] = layer_0[805] ^ layer_0[687]; 
    assign out[44] = layer_0[801] & layer_0[224]; 
    assign out[45] = layer_0[251] & layer_0[143]; 
    assign out[46] = ~layer_0[81]; 
    assign out[47] = ~(layer_0[1233] ^ layer_0[660]); 
    assign out[48] = layer_0[851] & layer_0[396]; 
    assign out[49] = layer_0[871] & ~layer_0[394]; 
    assign out[50] = ~layer_0[431] | (layer_0[449] & layer_0[431]); 
    assign out[51] = ~layer_0[653]; 
    assign out[52] = layer_0[1038] & ~layer_0[706]; 
    assign out[53] = layer_0[680]; 
    assign out[54] = layer_0[873] & ~layer_0[265]; 
    assign out[55] = ~(layer_0[1154] | layer_0[65]); 
    assign out[56] = ~layer_0[808] | (layer_0[6] & layer_0[808]); 
    assign out[57] = layer_0[275] & ~layer_0[725]; 
    assign out[58] = layer_0[642] | layer_0[710]; 
    assign out[59] = ~layer_0[1109]; 
    assign out[60] = layer_0[284]; 
    assign out[61] = layer_0[749] & ~layer_0[393]; 
    assign out[62] = layer_0[579] ^ layer_0[820]; 
    assign out[63] = ~layer_0[104]; 
    assign out[64] = layer_0[397] & ~layer_0[81]; 
    assign out[65] = ~(layer_0[68] ^ layer_0[476]); 
    assign out[66] = layer_0[660]; 
    assign out[67] = layer_0[559] ^ layer_0[506]; 
    assign out[68] = ~(layer_0[975] ^ layer_0[264]); 
    assign out[69] = layer_0[999] & layer_0[1049]; 
    assign out[70] = ~(layer_0[1085] ^ layer_0[949]); 
    assign out[71] = layer_0[341] ^ layer_0[488]; 
    assign out[72] = layer_0[966]; 
    assign out[73] = ~layer_0[588] | (layer_0[588] & layer_0[1204]); 
    assign out[74] = layer_0[1268] & ~layer_0[210]; 
    assign out[75] = layer_0[912] ^ layer_0[596]; 
    assign out[76] = layer_0[1025] & ~layer_0[297]; 
    assign out[77] = ~(layer_0[609] ^ layer_0[563]); 
    assign out[78] = ~layer_0[684]; 
    assign out[79] = layer_0[201] & layer_0[918]; 
    assign out[80] = ~(layer_0[38] & layer_0[60]); 
    assign out[81] = layer_0[517] | layer_0[312]; 
    assign out[82] = layer_0[492]; 
    assign out[83] = ~(layer_0[647] & layer_0[170]); 
    assign out[84] = layer_0[547]; 
    assign out[85] = ~layer_0[1226]; 
    assign out[86] = layer_0[566] & layer_0[770]; 
    assign out[87] = ~layer_0[1076]; 
    assign out[88] = ~(layer_0[1224] ^ layer_0[1257]); 
    assign out[89] = ~layer_0[1200] | (layer_0[1200] & layer_0[966]); 
    assign out[90] = layer_0[1257] & ~layer_0[464]; 
    assign out[91] = layer_0[341]; 
    assign out[92] = layer_0[995] & layer_0[1192]; 
    assign out[93] = layer_0[867]; 
    assign out[94] = layer_0[577] ^ layer_0[840]; 
    assign out[95] = layer_0[749] & ~layer_0[931]; 
    assign out[96] = ~(layer_0[550] ^ layer_0[54]); 
    assign out[97] = ~layer_0[499]; 
    assign out[98] = ~layer_0[636]; 
    assign out[99] = layer_0[1223] & layer_0[151]; 
    assign out[100] = layer_0[68] & layer_0[282]; 
    assign out[101] = layer_0[746] & ~layer_0[792]; 
    assign out[102] = layer_0[167] | layer_0[254]; 
    assign out[103] = ~layer_0[914]; 
    assign out[104] = ~(layer_0[1094] | layer_0[1225]); 
    assign out[105] = layer_0[100] ^ layer_0[1163]; 
    assign out[106] = ~(layer_0[1133] ^ layer_0[937]); 
    assign out[107] = layer_0[1104] ^ layer_0[1124]; 
    assign out[108] = ~layer_0[191] | (layer_0[572] & layer_0[191]); 
    assign out[109] = layer_0[908] & ~layer_0[655]; 
    assign out[110] = ~layer_0[819]; 
    assign out[111] = ~(layer_0[22] ^ layer_0[1050]); 
    assign out[112] = ~layer_0[931]; 
    assign out[113] = layer_0[481] & ~layer_0[331]; 
    assign out[114] = ~layer_0[508] | (layer_0[582] & layer_0[508]); 
    assign out[115] = ~(layer_0[1227] & layer_0[569]); 
    assign out[116] = layer_0[420]; 
    assign out[117] = ~(layer_0[1161] | layer_0[1127]); 
    assign out[118] = ~(layer_0[245] | layer_0[22]); 
    assign out[119] = layer_0[614]; 
    assign out[120] = layer_0[650] & ~layer_0[671]; 
    assign out[121] = layer_0[1140] & ~layer_0[63]; 
    assign out[122] = ~layer_0[983]; 
    assign out[123] = ~(layer_0[765] | layer_0[439]); 
    assign out[124] = ~(layer_0[162] | layer_0[243]); 
    assign out[125] = ~layer_0[60]; 
    assign out[126] = ~(layer_0[199] ^ layer_0[455]); 
    assign out[127] = ~layer_0[326] | (layer_0[1059] & layer_0[326]); 
    assign out[128] = ~(layer_0[1036] ^ layer_0[629]); 
    assign out[129] = layer_0[683] & ~layer_0[986]; 
    assign out[130] = ~layer_0[846]; 
    assign out[131] = ~layer_0[530]; 
    assign out[132] = layer_0[43]; 
    assign out[133] = layer_0[1263]; 
    assign out[134] = ~layer_0[1273] | (layer_0[1273] & layer_0[1009]); 
    assign out[135] = ~layer_0[133]; 
    assign out[136] = layer_0[1176]; 
    assign out[137] = layer_0[1165]; 
    assign out[138] = ~layer_0[1211]; 
    assign out[139] = ~layer_0[11] | (layer_0[797] & layer_0[11]); 
    assign out[140] = layer_0[936]; 
    assign out[141] = ~(layer_0[1192] ^ layer_0[1255]); 
    assign out[142] = ~layer_0[423] | (layer_0[423] & layer_0[1121]); 
    assign out[143] = ~(layer_0[223] ^ layer_0[555]); 
    assign out[144] = ~layer_0[693]; 
    assign out[145] = layer_0[1190]; 
    assign out[146] = layer_0[1183] & layer_0[395]; 
    assign out[147] = layer_0[988]; 
    assign out[148] = ~(layer_0[150] & layer_0[1182]); 
    assign out[149] = ~(layer_0[754] & layer_0[259]); 
    assign out[150] = layer_0[504] & ~layer_0[1249]; 
    assign out[151] = 1'b0; 
    assign out[152] = layer_0[634]; 
    assign out[153] = layer_0[489] ^ layer_0[750]; 
    assign out[154] = ~(layer_0[108] ^ layer_0[667]); 
    assign out[155] = layer_0[387] & ~layer_0[242]; 
    assign out[156] = ~(layer_0[1118] | layer_0[172]); 
    assign out[157] = layer_0[1120]; 
    assign out[158] = layer_0[1231]; 
    assign out[159] = layer_0[841]; 
    assign out[160] = ~(layer_0[595] ^ layer_0[1013]); 
    assign out[161] = ~(layer_0[1137] | layer_0[1258]); 
    assign out[162] = layer_0[1028] | layer_0[605]; 
    assign out[163] = ~(layer_0[695] ^ layer_0[1279]); 
    assign out[164] = layer_0[1073] & layer_0[257]; 
    assign out[165] = layer_0[711] ^ layer_0[778]; 
    assign out[166] = ~(layer_0[17] ^ layer_0[430]); 
    assign out[167] = ~(layer_0[944] ^ layer_0[489]); 
    assign out[168] = ~layer_0[89] | (layer_0[89] & layer_0[847]); 
    assign out[169] = layer_0[109] & ~layer_0[1161]; 
    assign out[170] = layer_0[573]; 
    assign out[171] = layer_0[1156] ^ layer_0[76]; 
    assign out[172] = ~(layer_0[1193] ^ layer_0[468]); 
    assign out[173] = layer_0[1240] & layer_0[187]; 
    assign out[174] = layer_0[1203] | layer_0[25]; 
    assign out[175] = layer_0[57]; 
    assign out[176] = layer_0[1154] ^ layer_0[866]; 
    assign out[177] = ~layer_0[985]; 
    assign out[178] = ~layer_0[20]; 
    assign out[179] = ~layer_0[1100]; 
    assign out[180] = layer_0[967] ^ layer_0[705]; 
    assign out[181] = layer_0[1016]; 
    assign out[182] = ~(layer_0[1081] ^ layer_0[514]); 
    assign out[183] = ~layer_0[523]; 
    assign out[184] = layer_0[880] ^ layer_0[678]; 
    assign out[185] = layer_0[509] ^ layer_0[1024]; 
    assign out[186] = ~layer_0[164]; 
    assign out[187] = layer_0[330] & layer_0[823]; 
    assign out[188] = ~(layer_0[1090] & layer_0[163]); 
    assign out[189] = layer_0[441] ^ layer_0[1160]; 
    assign out[190] = layer_0[373] & ~layer_0[457]; 
    assign out[191] = layer_0[1027] & ~layer_0[592]; 
    assign out[192] = ~layer_0[976] | (layer_0[368] & layer_0[976]); 
    assign out[193] = layer_0[500]; 
    assign out[194] = ~layer_0[190] | (layer_0[190] & layer_0[791]); 
    assign out[195] = layer_0[972] ^ layer_0[918]; 
    assign out[196] = ~layer_0[1033]; 
    assign out[197] = ~(layer_0[1117] ^ layer_0[292]); 
    assign out[198] = ~(layer_0[1093] ^ layer_0[469]); 
    assign out[199] = ~(layer_0[1223] ^ layer_0[610]); 
    assign out[200] = layer_0[704]; 
    assign out[201] = layer_0[442] ^ layer_0[436]; 
    assign out[202] = layer_0[703] ^ layer_0[501]; 
    assign out[203] = 1'b0; 
    assign out[204] = layer_0[359] & ~layer_0[515]; 
    assign out[205] = ~(layer_0[466] ^ layer_0[669]); 
    assign out[206] = ~(layer_0[1222] | layer_0[172]); 
    assign out[207] = ~(layer_0[298] | layer_0[180]); 
    assign out[208] = layer_0[1231] & ~layer_0[924]; 
    assign out[209] = layer_0[795]; 
    assign out[210] = ~(layer_0[244] ^ layer_0[405]); 
    assign out[211] = layer_0[676] & ~layer_0[283]; 
    assign out[212] = ~(layer_0[222] ^ layer_0[826]); 
    assign out[213] = layer_0[311] & ~layer_0[531]; 
    assign out[214] = layer_0[570] ^ layer_0[261]; 
    assign out[215] = ~(layer_0[277] ^ layer_0[376]); 
    assign out[216] = ~layer_0[941] | (layer_0[141] & layer_0[941]); 
    assign out[217] = ~(layer_0[555] ^ layer_0[148]); 
    assign out[218] = layer_0[24] & ~layer_0[408]; 
    assign out[219] = ~layer_0[325]; 
    assign out[220] = ~layer_0[354]; 
    assign out[221] = layer_0[847] & ~layer_0[635]; 
    assign out[222] = layer_0[152] & layer_0[1015]; 
    assign out[223] = layer_0[149] & ~layer_0[242]; 
    assign out[224] = ~(layer_0[945] | layer_0[753]); 
    assign out[225] = layer_0[411] & ~layer_0[998]; 
    assign out[226] = layer_0[468]; 
    assign out[227] = ~(layer_0[792] ^ layer_0[962]); 
    assign out[228] = ~(layer_0[1241] ^ layer_0[1077]); 
    assign out[229] = layer_0[659] ^ layer_0[321]; 
    assign out[230] = layer_0[827] ^ layer_0[375]; 
    assign out[231] = layer_0[971] & ~layer_0[1078]; 
    assign out[232] = layer_0[480] & ~layer_0[946]; 
    assign out[233] = layer_0[796]; 
    assign out[234] = ~(layer_0[729] ^ layer_0[1122]); 
    assign out[235] = layer_0[329]; 
    assign out[236] = layer_0[132] & ~layer_0[1063]; 
    assign out[237] = ~(layer_0[528] | layer_0[648]); 
    assign out[238] = layer_0[85] ^ layer_0[1032]; 
    assign out[239] = layer_0[795]; 
    assign out[240] = ~(layer_0[269] | layer_0[1137]); 
    assign out[241] = ~(layer_0[131] ^ layer_0[130]); 
    assign out[242] = layer_0[108] ^ layer_0[1214]; 
    assign out[243] = ~(layer_0[855] ^ layer_0[1044]); 
    assign out[244] = ~(layer_0[608] ^ layer_0[739]); 
    assign out[245] = layer_0[717] ^ layer_0[348]; 
    assign out[246] = ~(layer_0[727] | layer_0[5]); 
    assign out[247] = layer_0[665] ^ layer_0[688]; 
    assign out[248] = layer_0[206] ^ layer_0[602]; 
    assign out[249] = ~layer_0[1242]; 
    assign out[250] = ~layer_0[958] | (layer_0[550] & layer_0[958]); 
    assign out[251] = ~(layer_0[279] | layer_0[1098]); 
    assign out[252] = layer_0[318] ^ layer_0[917]; 
    assign out[253] = layer_0[77] & ~layer_0[457]; 
    assign out[254] = ~layer_0[640]; 
    assign out[255] = layer_0[843]; 
    assign out[256] = ~layer_0[861] | (layer_0[439] & layer_0[861]); 
    assign out[257] = layer_0[862] ^ layer_0[270]; 
    assign out[258] = layer_0[256]; 
    assign out[259] = layer_0[308] ^ layer_0[624]; 
    assign out[260] = layer_0[942]; 
    assign out[261] = ~(layer_0[565] ^ layer_0[895]); 
    assign out[262] = ~(layer_0[610] | layer_0[1100]); 
    assign out[263] = layer_0[557] ^ layer_0[799]; 
    assign out[264] = layer_0[7] | layer_0[356]; 
    assign out[265] = layer_0[725] & ~layer_0[1014]; 
    assign out[266] = layer_0[92] | layer_0[650]; 
    assign out[267] = layer_0[414] & layer_0[1019]; 
    assign out[268] = ~(layer_0[106] ^ layer_0[590]); 
    assign out[269] = ~(layer_0[406] ^ layer_0[235]); 
    assign out[270] = layer_0[851] ^ layer_0[1055]; 
    assign out[271] = ~layer_0[99] | (layer_0[252] & layer_0[99]); 
    assign out[272] = layer_0[628] ^ layer_0[788]; 
    assign out[273] = layer_0[1023] ^ layer_0[899]; 
    assign out[274] = layer_0[127]; 
    assign out[275] = ~(layer_0[1237] ^ layer_0[927]); 
    assign out[276] = layer_0[601]; 
    assign out[277] = ~layer_0[649]; 
    assign out[278] = ~(layer_0[91] ^ layer_0[572]); 
    assign out[279] = layer_0[930] & layer_0[916]; 
    assign out[280] = ~layer_0[154] | (layer_0[154] & layer_0[124]); 
    assign out[281] = layer_0[3] ^ layer_0[362]; 
    assign out[282] = ~layer_0[1113]; 
    assign out[283] = layer_0[1141] & ~layer_0[491]; 
    assign out[284] = layer_0[324]; 
    assign out[285] = layer_0[1217]; 
    assign out[286] = ~layer_0[970]; 
    assign out[287] = ~layer_0[516] | (layer_0[516] & layer_0[1083]); 
    assign out[288] = ~(layer_0[111] ^ layer_0[278]); 
    assign out[289] = ~(layer_0[593] ^ layer_0[1212]); 
    assign out[290] = layer_0[112] | layer_0[328]; 
    assign out[291] = layer_0[1078] ^ layer_0[692]; 
    assign out[292] = ~layer_0[1216]; 
    assign out[293] = layer_0[109] ^ layer_0[170]; 
    assign out[294] = ~(layer_0[475] ^ layer_0[784]); 
    assign out[295] = ~layer_0[456]; 
    assign out[296] = layer_0[574]; 
    assign out[297] = layer_0[928]; 
    assign out[298] = ~layer_0[1208]; 
    assign out[299] = layer_0[519] & ~layer_0[456]; 
    assign out[300] = ~(layer_0[1074] ^ layer_0[1091]); 
    assign out[301] = ~layer_0[560]; 
    assign out[302] = layer_0[839]; 
    assign out[303] = layer_0[904] | layer_0[327]; 
    assign out[304] = ~layer_0[754] | (layer_0[754] & layer_0[75]); 
    assign out[305] = layer_0[1211] ^ layer_0[906]; 
    assign out[306] = ~layer_0[959]; 
    assign out[307] = ~(layer_0[1261] & layer_0[346]); 
    assign out[308] = ~(layer_0[825] | layer_0[718]); 
    assign out[309] = ~layer_0[722] | (layer_0[500] & layer_0[722]); 
    assign out[310] = layer_0[1250] ^ layer_0[865]; 
    assign out[311] = ~layer_0[759]; 
    assign out[312] = layer_0[340]; 
    assign out[313] = ~(layer_0[1063] ^ layer_0[275]); 
    assign out[314] = layer_0[1159]; 
    assign out[315] = layer_0[1056] ^ layer_0[1067]; 
    assign out[316] = layer_0[91] & layer_0[490]; 
    assign out[317] = layer_0[234]; 
    assign out[318] = ~layer_0[342]; 
    assign out[319] = ~layer_0[458]; 
    assign out[320] = layer_0[295]; 
    assign out[321] = layer_0[599] ^ layer_0[1115]; 
    assign out[322] = ~layer_0[78]; 
    assign out[323] = layer_0[1226] & ~layer_0[556]; 
    assign out[324] = ~(layer_0[882] ^ layer_0[1130]); 
    assign out[325] = layer_0[878] ^ layer_0[454]; 
    assign out[326] = ~layer_0[1144] | (layer_0[1144] & layer_0[311]); 
    assign out[327] = layer_0[290]; 
    assign out[328] = layer_0[1037] ^ layer_0[767]; 
    assign out[329] = ~(layer_0[399] ^ layer_0[984]); 
    assign out[330] = ~layer_0[1196]; 
    assign out[331] = ~layer_0[144]; 
    assign out[332] = layer_0[306]; 
    assign out[333] = ~layer_0[189] | (layer_0[979] & layer_0[189]); 
    assign out[334] = ~(layer_0[357] ^ layer_0[71]); 
    assign out[335] = ~(layer_0[698] ^ layer_0[1004]); 
    assign out[336] = ~layer_0[1144] | (layer_0[811] & layer_0[1144]); 
    assign out[337] = layer_0[756]; 
    assign out[338] = layer_0[891]; 
    assign out[339] = ~(layer_0[615] | layer_0[887]); 
    assign out[340] = layer_0[1013] ^ layer_0[581]; 
    assign out[341] = layer_0[459]; 
    assign out[342] = ~layer_0[804]; 
    assign out[343] = layer_0[590] ^ layer_0[483]; 
    assign out[344] = ~layer_0[518] | (layer_0[897] & layer_0[518]); 
    assign out[345] = ~layer_0[198] | (layer_0[198] & layer_0[859]); 
    assign out[346] = layer_0[1251] ^ layer_0[471]; 
    assign out[347] = ~(layer_0[36] & layer_0[444]); 
    assign out[348] = layer_0[962]; 
    assign out[349] = ~layer_0[221]; 
    assign out[350] = layer_0[464] ^ layer_0[343]; 
    assign out[351] = layer_0[1000]; 
    assign out[352] = layer_0[318] & ~layer_0[452]; 
    assign out[353] = ~(layer_0[1] | layer_0[271]); 
    assign out[354] = layer_0[401] ^ layer_0[425]; 
    assign out[355] = layer_0[682] & layer_0[8]; 
    assign out[356] = ~layer_0[712]; 
    assign out[357] = ~(layer_0[314] ^ layer_0[415]); 
    assign out[358] = ~(layer_0[1124] ^ layer_0[619]); 
    assign out[359] = layer_0[222] | layer_0[216]; 
    assign out[360] = layer_0[312]; 
    assign out[361] = layer_0[674]; 
    assign out[362] = layer_0[447] & ~layer_0[789]; 
    assign out[363] = ~layer_0[309]; 
    assign out[364] = layer_0[961] & ~layer_0[1123]; 
    assign out[365] = ~layer_0[55] | (layer_0[6] & layer_0[55]); 
    assign out[366] = layer_0[916] & ~layer_0[330]; 
    assign out[367] = layer_0[933]; 
    assign out[368] = layer_0[130]; 
    assign out[369] = ~(layer_0[1072] ^ layer_0[1251]); 
    assign out[370] = ~(layer_0[478] & layer_0[834]); 
    assign out[371] = ~(layer_0[1075] ^ layer_0[424]); 
    assign out[372] = ~layer_0[970]; 
    assign out[373] = ~layer_0[591]; 
    assign out[374] = ~(layer_0[1170] | layer_0[745]); 
    assign out[375] = ~(layer_0[518] | layer_0[556]); 
    assign out[376] = layer_0[1064]; 
    assign out[377] = ~(layer_0[116] ^ layer_0[465]); 
    assign out[378] = layer_0[82] & layer_0[1000]; 
    assign out[379] = layer_0[186] & layer_0[447]; 
    assign out[380] = layer_0[1084] & ~layer_0[886]; 
    assign out[381] = layer_0[1006] & layer_0[485]; 
    assign out[382] = ~layer_0[87]; 
    assign out[383] = layer_0[365]; 
    assign out[384] = layer_0[1034] ^ layer_0[445]; 
    assign out[385] = layer_0[1209]; 
    assign out[386] = ~layer_0[121]; 
    assign out[387] = ~(layer_0[677] ^ layer_0[471]); 
    assign out[388] = ~layer_0[1229]; 
    assign out[389] = ~layer_0[817]; 
    assign out[390] = ~layer_0[522] | (layer_0[1225] & layer_0[522]); 
    assign out[391] = layer_0[320] | layer_0[757]; 
    assign out[392] = ~(layer_0[889] | layer_0[353]); 
    assign out[393] = ~layer_0[1220]; 
    assign out[394] = layer_0[594] ^ layer_0[380]; 
    assign out[395] = ~layer_0[536]; 
    assign out[396] = layer_0[115] ^ layer_0[418]; 
    assign out[397] = layer_0[16]; 
    assign out[398] = ~(layer_0[540] ^ layer_0[743]); 
    assign out[399] = layer_0[745]; 
    assign out[400] = ~layer_0[182]; 
    assign out[401] = layer_0[727] & ~layer_0[1051]; 
    assign out[402] = layer_0[248]; 
    assign out[403] = ~layer_0[463] | (layer_0[366] & layer_0[463]); 
    assign out[404] = ~(layer_0[882] ^ layer_0[1276]); 
    assign out[405] = layer_0[620]; 
    assign out[406] = layer_0[594]; 
    assign out[407] = ~layer_0[663]; 
    assign out[408] = layer_0[592]; 
    assign out[409] = ~(layer_0[1266] ^ layer_0[873]); 
    assign out[410] = ~(layer_0[626] ^ layer_0[51]); 
    assign out[411] = layer_0[1069]; 
    assign out[412] = ~layer_0[934]; 
    assign out[413] = layer_0[371]; 
    assign out[414] = layer_0[186] & ~layer_0[1193]; 
    assign out[415] = layer_0[950]; 
    assign out[416] = ~layer_0[229]; 
    assign out[417] = ~(layer_0[923] | layer_0[1019]); 
    assign out[418] = ~(layer_0[1004] ^ layer_0[90]); 
    assign out[419] = layer_0[965] & ~layer_0[1097]; 
    assign out[420] = layer_0[542] ^ layer_0[412]; 
    assign out[421] = layer_0[676]; 
    assign out[422] = ~layer_0[14]; 
    assign out[423] = ~(layer_0[1041] & layer_0[568]); 
    assign out[424] = ~(layer_0[233] & layer_0[711]); 
    assign out[425] = ~layer_0[1048]; 
    assign out[426] = ~layer_0[104]; 
    assign out[427] = ~(layer_0[443] ^ layer_0[965]); 
    assign out[428] = layer_0[192] & layer_0[709]; 
    assign out[429] = ~(layer_0[757] ^ layer_0[760]); 
    assign out[430] = layer_0[937] & ~layer_0[1140]; 
    assign out[431] = ~(layer_0[1082] ^ layer_0[781]); 
    assign out[432] = ~layer_0[260]; 
    assign out[433] = layer_0[744] & ~layer_0[580]; 
    assign out[434] = layer_0[1029]; 
    assign out[435] = layer_0[340]; 
    assign out[436] = ~layer_0[36]; 
    assign out[437] = ~layer_0[579]; 
    assign out[438] = ~layer_0[1169]; 
    assign out[439] = layer_0[748]; 
    assign out[440] = layer_0[392] ^ layer_0[1219]; 
    assign out[441] = ~(layer_0[443] ^ layer_0[493]); 
    assign out[442] = layer_0[460] ^ layer_0[159]; 
    assign out[443] = layer_0[147] & ~layer_0[604]; 
    assign out[444] = layer_0[198] ^ layer_0[440]; 
    assign out[445] = ~layer_0[503]; 
    assign out[446] = layer_0[118]; 
    assign out[447] = layer_0[1275] ^ layer_0[779]; 
    assign out[448] = layer_0[389] ^ layer_0[42]; 
    assign out[449] = ~(layer_0[929] ^ layer_0[977]); 
    assign out[450] = layer_0[808] ^ layer_0[677]; 
    assign out[451] = ~layer_0[301]; 
    assign out[452] = ~(layer_0[482] ^ layer_0[1246]); 
    assign out[453] = layer_0[204] & ~layer_0[557]; 
    assign out[454] = ~layer_0[73]; 
    assign out[455] = layer_0[241] ^ layer_0[801]; 
    assign out[456] = layer_0[600] ^ layer_0[770]; 
    assign out[457] = layer_0[490] & ~layer_0[1020]; 
    assign out[458] = ~(layer_0[250] ^ layer_0[1239]); 
    assign out[459] = ~layer_0[503] | (layer_0[595] & layer_0[503]); 
    assign out[460] = ~(layer_0[136] ^ layer_0[865]); 
    assign out[461] = ~(layer_0[641] ^ layer_0[369]); 
    assign out[462] = ~layer_0[874] | (layer_0[67] & layer_0[874]); 
    assign out[463] = layer_0[123]; 
    assign out[464] = ~layer_0[23]; 
    assign out[465] = layer_0[317] | layer_0[332]; 
    assign out[466] = ~layer_0[1075]; 
    assign out[467] = layer_0[621] ^ layer_0[304]; 
    assign out[468] = layer_0[672]; 
    assign out[469] = layer_0[831] & layer_0[70]; 
    assign out[470] = layer_0[696]; 
    assign out[471] = layer_0[583] & ~layer_0[453]; 
    assign out[472] = layer_0[763]; 
    assign out[473] = ~(layer_0[1172] & layer_0[343]); 
    assign out[474] = layer_0[1207] | layer_0[52]; 
    assign out[475] = layer_0[1053] | layer_0[136]; 
    assign out[476] = ~(layer_0[97] ^ layer_0[1068]); 
    assign out[477] = layer_0[658] ^ layer_0[157]; 
    assign out[478] = ~layer_0[467]; 
    assign out[479] = layer_0[517] ^ layer_0[751]; 
    assign out[480] = layer_0[472] & ~layer_0[746]; 
    assign out[481] = ~layer_0[1277] | (layer_0[900] & layer_0[1277]); 
    assign out[482] = layer_0[32] | layer_0[1042]; 
    assign out[483] = layer_0[448]; 
    assign out[484] = layer_0[891]; 
    assign out[485] = ~layer_0[177]; 
    assign out[486] = ~layer_0[446]; 
    assign out[487] = layer_0[56] ^ layer_0[758]; 
    assign out[488] = layer_0[295] ^ layer_0[863]; 
    assign out[489] = layer_0[352]; 
    assign out[490] = layer_0[128] & ~layer_0[157]; 
    assign out[491] = layer_0[841] ^ layer_0[686]; 
    assign out[492] = layer_0[477] & ~layer_0[384]; 
    assign out[493] = ~(layer_0[675] ^ layer_0[189]); 
    assign out[494] = layer_0[681]; 
    assign out[495] = ~(layer_0[744] ^ layer_0[347]); 
    assign out[496] = ~layer_0[597]; 
    assign out[497] = layer_0[734] & ~layer_0[281]; 
    assign out[498] = layer_0[145]; 
    assign out[499] = ~(layer_0[302] ^ layer_0[993]); 
    assign out[500] = ~(layer_0[215] ^ layer_0[619]); 
    assign out[501] = layer_0[575]; 
    assign out[502] = ~(layer_0[376] ^ layer_0[513]); 
    assign out[503] = ~layer_0[783] | (layer_0[783] & layer_0[200]); 
    assign out[504] = ~layer_0[876]; 
    assign out[505] = ~(layer_0[765] ^ layer_0[812]); 
    assign out[506] = layer_0[967] ^ layer_0[285]; 
    assign out[507] = ~(layer_0[1127] ^ layer_0[992]); 
    assign out[508] = ~layer_0[1195]; 
    assign out[509] = layer_0[1027] & ~layer_0[422]; 
    assign out[510] = ~(layer_0[240] | layer_0[424]); 
    assign out[511] = ~(layer_0[327] ^ layer_0[726]); 
    assign out[512] = ~layer_0[774]; 
    assign out[513] = layer_0[607] ^ layer_0[180]; 
    assign out[514] = layer_0[989] & layer_0[662]; 
    assign out[515] = ~layer_0[694]; 
    assign out[516] = ~(layer_0[762] ^ layer_0[992]); 
    assign out[517] = layer_0[301]; 
    assign out[518] = layer_0[264]; 
    assign out[519] = layer_0[528]; 
    assign out[520] = ~layer_0[1001]; 
    assign out[521] = layer_0[135] & ~layer_0[310]; 
    assign out[522] = ~(layer_0[1139] ^ layer_0[1079]); 
    assign out[523] = layer_0[263] & layer_0[1185]; 
    assign out[524] = layer_0[558] ^ layer_0[117]; 
    assign out[525] = layer_0[329] & layer_0[668]; 
    assign out[526] = ~(layer_0[630] | layer_0[4]); 
    assign out[527] = layer_0[1112]; 
    assign out[528] = layer_0[858] ^ layer_0[44]; 
    assign out[529] = layer_0[544] ^ layer_0[1245]; 
    assign out[530] = ~layer_0[409]; 
    assign out[531] = ~layer_0[1267] | (layer_0[1267] & layer_0[334]); 
    assign out[532] = ~layer_0[266]; 
    assign out[533] = layer_0[1003] & ~layer_0[601]; 
    assign out[534] = layer_0[165] ^ layer_0[505]; 
    assign out[535] = layer_0[1050] ^ layer_0[433]; 
    assign out[536] = ~(layer_0[761] ^ layer_0[545]); 
    assign out[537] = ~(layer_0[268] | layer_0[80]); 
    assign out[538] = layer_0[1048] & layer_0[404]; 
    assign out[539] = layer_0[412]; 
    assign out[540] = layer_0[360]; 
    assign out[541] = layer_0[889]; 
    assign out[542] = ~(layer_0[955] | layer_0[645]); 
    assign out[543] = ~(layer_0[1156] ^ layer_0[1155]); 
    assign out[544] = ~layer_0[350]; 
    assign out[545] = layer_0[1159] ^ layer_0[997]; 
    assign out[546] = layer_0[495]; 
    assign out[547] = ~(layer_0[1134] | layer_0[854]); 
    assign out[548] = layer_0[887]; 
    assign out[549] = ~layer_0[338]; 
    assign out[550] = layer_0[44] ^ layer_0[1175]; 
    assign out[551] = layer_0[816] & ~layer_0[633]; 
    assign out[552] = layer_0[960] | layer_0[1178]; 
    assign out[553] = layer_0[1086] ^ layer_0[999]; 
    assign out[554] = ~(layer_0[142] | layer_0[736]); 
    assign out[555] = ~layer_0[1117] | (layer_0[143] & layer_0[1117]); 
    assign out[556] = ~(layer_0[943] ^ layer_0[1273]); 
    assign out[557] = layer_0[892]; 
    assign out[558] = layer_0[185] & ~layer_0[864]; 
    assign out[559] = layer_0[625] ^ layer_0[713]; 
    assign out[560] = layer_0[194]; 
    assign out[561] = ~(layer_0[521] ^ layer_0[1057]); 
    assign out[562] = ~(layer_0[996] ^ layer_0[441]); 
    assign out[563] = layer_0[1196] ^ layer_0[357]; 
    assign out[564] = layer_0[19]; 
    assign out[565] = ~layer_0[101]; 
    assign out[566] = ~(layer_0[42] ^ layer_0[298]); 
    assign out[567] = ~layer_0[1164]; 
    assign out[568] = ~layer_0[35] | (layer_0[207] & layer_0[35]); 
    assign out[569] = ~(layer_0[656] ^ layer_0[37]); 
    assign out[570] = layer_0[853] & ~layer_0[569]; 
    assign out[571] = ~layer_0[1028]; 
    assign out[572] = ~layer_0[1207]; 
    assign out[573] = ~layer_0[20]; 
    assign out[574] = ~layer_0[274]; 
    assign out[575] = ~(layer_0[781] ^ layer_0[1017]); 
    assign out[576] = layer_0[1044] | layer_0[1150]; 
    assign out[577] = layer_0[207] & ~layer_0[296]; 
    assign out[578] = ~layer_0[455]; 
    assign out[579] = layer_0[74] & layer_0[102]; 
    assign out[580] = layer_0[273] & ~layer_0[573]; 
    assign out[581] = ~(layer_0[105] ^ layer_0[491]); 
    assign out[582] = layer_0[828] & layer_0[349]; 
    assign out[583] = layer_0[1046] ^ layer_0[648]; 
    assign out[584] = ~(layer_0[605] ^ layer_0[1208]); 
    assign out[585] = ~(layer_0[1015] ^ layer_0[1254]); 
    assign out[586] = ~(layer_0[1052] | layer_0[155]); 
    assign out[587] = ~(layer_0[673] ^ layer_0[654]); 
    assign out[588] = layer_0[525] | layer_0[286]; 
    assign out[589] = ~layer_0[98]; 
    assign out[590] = ~layer_0[307]; 
    assign out[591] = ~(layer_0[618] ^ layer_0[50]); 
    assign out[592] = ~layer_0[1165]; 
    assign out[593] = layer_0[470]; 
    assign out[594] = ~(layer_0[1253] ^ layer_0[849]); 
    assign out[595] = ~layer_0[1069]; 
    assign out[596] = ~(layer_0[220] ^ layer_0[577]); 
    assign out[597] = ~layer_0[418]; 
    assign out[598] = layer_0[1201] & layer_0[358]; 
    assign out[599] = layer_0[599] ^ layer_0[432]; 
    assign out[600] = layer_0[718]; 
    assign out[601] = layer_0[901] & ~layer_0[616]; 
    assign out[602] = ~(layer_0[1179] ^ layer_0[299]); 
    assign out[603] = ~layer_0[1052] | (layer_0[1052] & layer_0[1119]); 
    assign out[604] = ~(layer_0[979] ^ layer_0[731]); 
    assign out[605] = ~(layer_0[768] ^ layer_0[567]); 
    assign out[606] = layer_0[1126]; 
    assign out[607] = ~layer_0[370]; 
    assign out[608] = ~(layer_0[332] ^ layer_0[827]); 
    assign out[609] = layer_0[476] ^ layer_0[524]; 
    assign out[610] = layer_0[362] ^ layer_0[171]; 
    assign out[611] = ~layer_0[165] | (layer_0[165] & layer_0[334]); 
    assign out[612] = ~(layer_0[208] & layer_0[1190]); 
    assign out[613] = layer_0[446] & ~layer_0[1274]; 
    assign out[614] = layer_0[939] ^ layer_0[836]; 
    assign out[615] = layer_0[1256] & ~layer_0[790]; 
    assign out[616] = ~layer_0[533]; 
    assign out[617] = ~layer_0[649]; 
    assign out[618] = layer_0[391] ^ layer_0[585]; 
    assign out[619] = ~(layer_0[687] & layer_0[375]); 
    assign out[620] = layer_0[294] ^ layer_0[561]; 
    assign out[621] = layer_0[902] ^ layer_0[606]; 
    assign out[622] = ~(layer_0[775] ^ layer_0[838]); 
    assign out[623] = layer_0[842] & layer_0[54]; 
    assign out[624] = ~layer_0[630]; 
    assign out[625] = layer_0[1173] & layer_0[1030]; 
    assign out[626] = layer_0[773] ^ layer_0[474]; 
    assign out[627] = ~layer_0[378] | (layer_0[171] & layer_0[378]); 
    assign out[628] = layer_0[299] ^ layer_0[213]; 
    assign out[629] = layer_0[493] ^ layer_0[982]; 
    assign out[630] = layer_0[802] ^ layer_0[348]; 
    assign out[631] = layer_0[959] ^ layer_0[342]; 
    assign out[632] = layer_0[829] & layer_0[1098]; 
    assign out[633] = ~(layer_0[1215] ^ layer_0[139]); 
    assign out[634] = ~layer_0[657] | (layer_0[133] & layer_0[657]); 
    assign out[635] = layer_0[1088] ^ layer_0[276]; 
    assign out[636] = ~layer_0[64]; 
    assign out[637] = layer_0[1158]; 
    assign out[638] = ~(layer_0[141] & layer_0[403]); 
    assign out[639] = layer_0[1061] ^ layer_0[688]; 
    assign out[640] = layer_0[382]; 
    assign out[641] = ~(layer_0[850] & layer_0[1073]); 
    assign out[642] = layer_0[88] & ~layer_0[584]; 
    assign out[643] = layer_0[1108] ^ layer_0[643]; 
    assign out[644] = layer_0[325]; 
    assign out[645] = layer_0[1263] ^ layer_0[670]; 
    assign out[646] = layer_0[1090] ^ layer_0[939]; 
    assign out[647] = ~(layer_0[886] ^ layer_0[1129]); 
    assign out[648] = layer_0[609] ^ layer_0[1011]; 
    assign out[649] = ~(layer_0[303] ^ layer_0[1182]); 
    assign out[650] = layer_0[1242]; 
    assign out[651] = layer_0[379] ^ layer_0[1120]; 
    assign out[652] = layer_0[1095]; 
    assign out[653] = ~(layer_0[344] ^ layer_0[444]); 
    assign out[654] = ~layer_0[627] | (layer_0[735] & layer_0[627]); 
    assign out[655] = layer_0[220] ^ layer_0[537]; 
    assign out[656] = ~layer_0[1162]; 
    assign out[657] = ~layer_0[707]; 
    assign out[658] = ~layer_0[769]; 
    assign out[659] = ~(layer_0[640] & layer_0[1053]); 
    assign out[660] = ~layer_0[323] | (layer_0[323] & layer_0[715]); 
    assign out[661] = layer_0[848]; 
    assign out[662] = ~layer_0[1057] | (layer_0[1057] & layer_0[185]); 
    assign out[663] = ~(layer_0[1244] ^ layer_0[708]); 
    assign out[664] = ~(layer_0[818] | layer_0[272]); 
    assign out[665] = ~layer_0[859] | (layer_0[859] & layer_0[113]); 
    assign out[666] = layer_0[739] & ~layer_0[645]; 
    assign out[667] = ~(layer_0[282] ^ layer_0[1094]); 
    assign out[668] = ~layer_0[596]; 
    assign out[669] = ~layer_0[74] | (layer_0[146] & layer_0[74]); 
    assign out[670] = ~(layer_0[836] ^ layer_0[497]); 
    assign out[671] = layer_0[520]; 
    assign out[672] = layer_0[868]; 
    assign out[673] = ~layer_0[1009]; 
    assign out[674] = layer_0[532] ^ layer_0[230]; 
    assign out[675] = layer_0[668]; 
    assign out[676] = ~layer_0[831] | (layer_0[169] & layer_0[831]); 
    assign out[677] = layer_0[719] ^ layer_0[685]; 
    assign out[678] = layer_0[1] | layer_0[17]; 
    assign out[679] = ~(layer_0[671] ^ layer_0[237]); 
    assign out[680] = layer_0[664]; 
    assign out[681] = ~layer_0[885]; 
    assign out[682] = layer_0[1107] ^ layer_0[1089]; 
    assign out[683] = ~layer_0[179] | (layer_0[216] & layer_0[179]); 
    assign out[684] = layer_0[534]; 
    assign out[685] = ~(layer_0[661] & layer_0[1184]); 
    assign out[686] = layer_0[637]; 
    assign out[687] = layer_0[256] ^ layer_0[1197]; 
    assign out[688] = layer_0[173]; 
    assign out[689] = ~(layer_0[13] | layer_0[1247]); 
    assign out[690] = ~(layer_0[627] | layer_0[358]); 
    assign out[691] = layer_0[465] ^ layer_0[1007]; 
    assign out[692] = ~layer_0[1221] | (layer_0[1221] & layer_0[789]); 
    assign out[693] = ~(layer_0[333] ^ layer_0[112]); 
    assign out[694] = layer_0[697] ^ layer_0[137]; 
    assign out[695] = ~(layer_0[1136] & layer_0[608]); 
    assign out[696] = layer_0[613] ^ layer_0[249]; 
    assign out[697] = layer_0[353] ^ layer_0[237]; 
    assign out[698] = ~layer_0[265] | (layer_0[435] & layer_0[265]); 
    assign out[699] = ~layer_0[1217]; 
    assign out[700] = layer_0[915] ^ layer_0[414]; 
    assign out[701] = ~(layer_0[913] ^ layer_0[552]); 
    assign out[702] = ~layer_0[584]; 
    assign out[703] = layer_0[1095] | layer_0[197]; 
    assign out[704] = ~(layer_0[402] ^ layer_0[763]); 
    assign out[705] = ~(layer_0[434] ^ layer_0[230]); 
    assign out[706] = ~layer_0[885]; 
    assign out[707] = ~(layer_0[954] ^ layer_0[1139]); 
    assign out[708] = layer_0[238] ^ layer_0[663]; 
    assign out[709] = layer_0[666]; 
    assign out[710] = layer_0[178] & ~layer_0[856]; 
    assign out[711] = layer_0[307]; 
    assign out[712] = layer_0[893] & ~layer_0[46]; 
    assign out[713] = layer_0[777] | layer_0[1056]; 
    assign out[714] = layer_0[691] | layer_0[219]; 
    assign out[715] = layer_0[1243]; 
    assign out[716] = ~layer_0[138] | (layer_0[138] & layer_0[951]); 
    assign out[717] = layer_0[482] ^ layer_0[1096]; 
    assign out[718] = layer_0[485] ^ layer_0[624]; 
    assign out[719] = ~(layer_0[1205] ^ layer_0[786]); 
    assign out[720] = ~(layer_0[898] ^ layer_0[580]); 
    assign out[721] = layer_0[860] & layer_0[512]; 
    assign out[722] = layer_0[602]; 
    assign out[723] = ~layer_0[1174]; 
    assign out[724] = ~layer_0[850] | (layer_0[466] & layer_0[850]); 
    assign out[725] = layer_0[783]; 
    assign out[726] = layer_0[629] | layer_0[907]; 
    assign out[727] = layer_0[554] ^ layer_0[206]; 
    assign out[728] = layer_0[253]; 
    assign out[729] = layer_0[696]; 
    assign out[730] = ~layer_0[84] | (layer_0[84] & layer_0[29]); 
    assign out[731] = ~(layer_0[344] ^ layer_0[492]); 
    assign out[732] = ~layer_0[1084]; 
    assign out[733] = layer_0[119] | layer_0[1167]; 
    assign out[734] = ~(layer_0[53] ^ layer_0[335]); 
    assign out[735] = layer_0[620]; 
    assign out[736] = layer_0[824]; 
    assign out[737] = ~(layer_0[1022] ^ layer_0[720]); 
    assign out[738] = layer_0[587]; 
    assign out[739] = ~(layer_0[126] ^ layer_0[372]); 
    assign out[740] = layer_0[614]; 
    assign out[741] = ~(layer_0[26] ^ layer_0[913]); 
    assign out[742] = ~layer_0[707]; 
    assign out[743] = ~(layer_0[478] & layer_0[527]); 
    assign out[744] = layer_0[777] ^ layer_0[23]; 
    assign out[745] = ~(layer_0[879] ^ layer_0[365]); 
    assign out[746] = layer_0[274] & layer_0[35]; 
    assign out[747] = ~(layer_0[541] ^ layer_0[63]); 
    assign out[748] = ~(layer_0[844] & layer_0[578]); 
    assign out[749] = ~layer_0[28] | (layer_0[28] & layer_0[1093]); 
    assign out[750] = ~layer_0[632]; 
    assign out[751] = ~layer_0[1188]; 
    assign out[752] = ~(layer_0[1204] ^ layer_0[469]); 
    assign out[753] = layer_0[549] ^ layer_0[434]; 
    assign out[754] = ~(layer_0[521] ^ layer_0[715]); 
    assign out[755] = ~(layer_0[184] ^ layer_0[737]); 
    assign out[756] = layer_0[395]; 
    assign out[757] = ~layer_0[486] | (layer_0[486] & layer_0[58]); 
    assign out[758] = ~layer_0[802]; 
    assign out[759] = ~layer_0[538] | (layer_0[753] & layer_0[538]); 
    assign out[760] = layer_0[1276]; 
    assign out[761] = layer_0[413] ^ layer_0[287]; 
    assign out[762] = layer_0[438]; 
    assign out[763] = layer_0[1131] | layer_0[392]; 
    assign out[764] = ~(layer_0[911] | layer_0[935]); 
    assign out[765] = layer_0[87] & layer_0[1232]; 
    assign out[766] = layer_0[1006]; 
    assign out[767] = ~layer_0[31]; 
    assign out[768] = ~(layer_0[371] | layer_0[226]); 
    assign out[769] = ~(layer_0[1210] | layer_0[320]); 
    assign out[770] = layer_0[270] & layer_0[208]; 
    assign out[771] = ~layer_0[251]; 
    assign out[772] = ~layer_0[659]; 
    assign out[773] = layer_0[654] & ~layer_0[429]; 
    assign out[774] = ~(layer_0[1141] & layer_0[582]); 
    assign out[775] = layer_0[558]; 
    assign out[776] = ~(layer_0[733] | layer_0[656]); 
    assign out[777] = ~layer_0[898] | (layer_0[898] & layer_0[66]); 
    assign out[778] = layer_0[946]; 
    assign out[779] = layer_0[419] | layer_0[742]; 
    assign out[780] = layer_0[904] & ~layer_0[604]; 
    assign out[781] = ~layer_0[1018] | (layer_0[1018] & layer_0[615]); 
    assign out[782] = layer_0[494] ^ layer_0[1186]; 
    assign out[783] = layer_0[310] ^ layer_0[1163]; 
    assign out[784] = layer_0[1023] & ~layer_0[1022]; 
    assign out[785] = ~(layer_0[79] ^ layer_0[8]); 
    assign out[786] = ~layer_0[364]; 
    assign out[787] = ~(layer_0[2] | layer_0[161]); 
    assign out[788] = layer_0[1003] & ~layer_0[1108]; 
    assign out[789] = layer_0[473]; 
    assign out[790] = layer_0[93] ^ layer_0[994]; 
    assign out[791] = layer_0[700] & layer_0[987]; 
    assign out[792] = layer_0[1102] & ~layer_0[1143]; 
    assign out[793] = layer_0[1110] ^ layer_0[778]; 
    assign out[794] = ~(layer_0[1210] & layer_0[147]); 
    assign out[795] = ~(layer_0[719] ^ layer_0[1184]); 
    assign out[796] = ~(layer_0[58] ^ layer_0[597]); 
    assign out[797] = layer_0[515] & layer_0[690]; 
    assign out[798] = layer_0[1147]; 
    assign out[799] = layer_0[583] & ~layer_0[1176]; 
    assign out[800] = layer_0[1271] & ~layer_0[235]; 
    assign out[801] = ~(layer_0[636] | layer_0[978]); 
    assign out[802] = layer_0[1220] & ~layer_0[135]; 
    assign out[803] = ~(layer_0[603] ^ layer_0[787]); 
    assign out[804] = layer_0[948] ^ layer_0[586]; 
    assign out[805] = ~(layer_0[132] ^ layer_0[1185]); 
    assign out[806] = layer_0[1214] | layer_0[1240]; 
    assign out[807] = layer_0[1195] & ~layer_0[1008]; 
    assign out[808] = layer_0[643] & ~layer_0[673]; 
    assign out[809] = ~(layer_0[984] & layer_0[911]); 
    assign out[810] = ~(layer_0[723] ^ layer_0[27]); 
    assign out[811] = layer_0[1026] & layer_0[945]; 
    assign out[812] = layer_0[285] & ~layer_0[1166]; 
    assign out[813] = ~layer_0[1010]; 
    assign out[814] = ~layer_0[138]; 
    assign out[815] = layer_0[1238]; 
    assign out[816] = layer_0[148]; 
    assign out[817] = layer_0[938] & layer_0[352]; 
    assign out[818] = layer_0[142] ^ layer_0[864]; 
    assign out[819] = ~layer_0[822] | (layer_0[822] & layer_0[869]); 
    assign out[820] = layer_0[1262] ^ layer_0[575]; 
    assign out[821] = ~layer_0[168]; 
    assign out[822] = layer_0[972] & ~layer_0[487]; 
    assign out[823] = ~layer_0[477]; 
    assign out[824] = layer_0[24] & ~layer_0[638]; 
    assign out[825] = layer_0[1148]; 
    assign out[826] = layer_0[987] & ~layer_0[1034]; 
    assign out[827] = ~layer_0[423]; 
    assign out[828] = layer_0[662] & ~layer_0[1241]; 
    assign out[829] = layer_0[695] ^ layer_0[1105]; 
    assign out[830] = layer_0[1103] & ~layer_0[564]; 
    assign out[831] = ~layer_0[46] | (layer_0[355] & layer_0[46]); 
    assign out[832] = ~(layer_0[367] ^ layer_0[903]); 
    assign out[833] = layer_0[345] ^ layer_0[1115]; 
    assign out[834] = ~(layer_0[552] ^ layer_0[41]); 
    assign out[835] = ~(layer_0[1092] ^ layer_0[646]); 
    assign out[836] = layer_0[800]; 
    assign out[837] = ~(layer_0[1259] ^ layer_0[699]); 
    assign out[838] = ~layer_0[31]; 
    assign out[839] = ~(layer_0[733] | layer_0[1101]); 
    assign out[840] = ~layer_0[546] | (layer_0[498] & layer_0[546]); 
    assign out[841] = ~(layer_0[123] | layer_0[1077]); 
    assign out[842] = layer_0[807]; 
    assign out[843] = layer_0[1002] & ~layer_0[1202]; 
    assign out[844] = layer_0[1114] ^ layer_0[101]; 
    assign out[845] = ~layer_0[271]; 
    assign out[846] = ~(layer_0[764] ^ layer_0[11]); 
    assign out[847] = layer_0[571] ^ layer_0[701]; 
    assign out[848] = layer_0[335]; 
    assign out[849] = ~layer_0[899] | (layer_0[111] & layer_0[899]); 
    assign out[850] = layer_0[986]; 
    assign out[851] = ~layer_0[153]; 
    assign out[852] = layer_0[1135] ^ layer_0[1152]; 
    assign out[853] = layer_0[1168] & ~layer_0[798]; 
    assign out[854] = ~(layer_0[1261] | layer_0[1110]); 
    assign out[855] = layer_0[973] & ~layer_0[914]; 
    assign out[856] = ~(layer_0[566] ^ layer_0[807]); 
    assign out[857] = ~layer_0[1065] | (layer_0[88] & layer_0[1065]); 
    assign out[858] = layer_0[639]; 
    assign out[859] = layer_0[647] & ~layer_0[787]; 
    assign out[860] = ~(layer_0[724] ^ layer_0[415]); 
    assign out[861] = ~(layer_0[1131] ^ layer_0[1187]); 
    assign out[862] = ~layer_0[644] | (layer_0[1123] & layer_0[644]); 
    assign out[863] = layer_0[845] & layer_0[871]; 
    assign out[864] = ~(layer_0[1157] & layer_0[883]); 
    assign out[865] = ~layer_0[304] | (layer_0[1262] & layer_0[304]); 
    assign out[866] = ~layer_0[861]; 
    assign out[867] = ~(layer_0[511] ^ layer_0[153]); 
    assign out[868] = layer_0[1054] & layer_0[1002]; 
    assign out[869] = layer_0[724] | layer_0[526]; 
    assign out[870] = ~(layer_0[598] ^ layer_0[78]); 
    assign out[871] = layer_0[1199] & ~layer_0[253]; 
    assign out[872] = layer_0[462] & layer_0[45]; 
    assign out[873] = ~layer_0[969]; 
    assign out[874] = ~layer_0[303]; 
    assign out[875] = ~(layer_0[323] ^ layer_0[722]); 
    assign out[876] = layer_0[261]; 
    assign out[877] = ~layer_0[562]; 
    assign out[878] = ~layer_0[1191]; 
    assign out[879] = layer_0[209]; 
    assign out[880] = layer_0[1007] & ~layer_0[239]; 
    assign out[881] = ~(layer_0[679] ^ layer_0[1275]); 
    assign out[882] = layer_0[337] & ~layer_0[928]; 
    assign out[883] = ~(layer_0[990] | layer_0[156]); 
    assign out[884] = ~layer_0[313]; 
    assign out[885] = ~(layer_0[1200] ^ layer_0[246]); 
    assign out[886] = layer_0[666]; 
    assign out[887] = ~layer_0[283] | (layer_0[926] & layer_0[283]); 
    assign out[888] = ~layer_0[1246]; 
    assign out[889] = ~layer_0[721]; 
    assign out[890] = ~layer_0[177]; 
    assign out[891] = ~(layer_0[1151] ^ layer_0[445]); 
    assign out[892] = ~layer_0[1058] | (layer_0[998] & layer_0[1058]); 
    assign out[893] = layer_0[1142] & ~layer_0[935]; 
    assign out[894] = ~(layer_0[798] | layer_0[679]); 
    assign out[895] = ~(layer_0[824] ^ layer_0[1212]); 
    assign out[896] = ~layer_0[675]; 
    assign out[897] = ~layer_0[879]; 
    assign out[898] = ~(layer_0[427] ^ layer_0[174]); 
    assign out[899] = layer_0[387] ^ layer_0[398]; 
    assign out[900] = layer_0[115] | layer_0[291]; 
    assign out[901] = ~(layer_0[67] ^ layer_0[922]); 
    assign out[902] = ~layer_0[1062]; 
    assign out[903] = layer_0[461] | layer_0[229]; 
    assign out[904] = ~layer_0[1158]; 
    assign out[905] = ~layer_0[288] | (layer_0[288] & layer_0[199]); 
    assign out[906] = layer_0[337] ^ layer_0[350]; 
    assign out[907] = ~layer_0[912]; 
    assign out[908] = ~layer_0[842] | (layer_0[842] & layer_0[66]); 
    assign out[909] = ~(layer_0[113] ^ layer_0[62]); 
    assign out[910] = ~(layer_0[80] ^ layer_0[117]); 
    assign out[911] = layer_0[203] ^ layer_0[225]; 
    assign out[912] = layer_0[1080] & layer_0[94]; 
    assign out[913] = layer_0[717]; 
    assign out[914] = ~(layer_0[10] | layer_0[699]); 
    assign out[915] = layer_0[883] & ~layer_0[33]; 
    assign out[916] = layer_0[835]; 
    assign out[917] = ~(layer_0[728] | layer_0[249]); 
    assign out[918] = ~(layer_0[227] ^ layer_0[603]); 
    assign out[919] = layer_0[409]; 
    assign out[920] = ~layer_0[682]; 
    assign out[921] = layer_0[564]; 
    assign out[922] = ~layer_0[48]; 
    assign out[923] = layer_0[920] & ~layer_0[755]; 
    assign out[924] = layer_0[1157] | layer_0[145]; 
    assign out[925] = layer_0[416] & layer_0[1082]; 
    assign out[926] = layer_0[723] ^ layer_0[12]; 
    assign out[927] = ~(layer_0[941] | layer_0[160]); 
    assign out[928] = layer_0[168] & ~layer_0[638]; 
    assign out[929] = ~(layer_0[706] ^ layer_0[821]); 
    assign out[930] = layer_0[1235] ^ layer_0[289]; 
    assign out[931] = layer_0[774]; 
    assign out[932] = layer_0[785] ^ layer_0[70]; 
    assign out[933] = ~(layer_0[1248] ^ layer_0[194]); 
    assign out[934] = ~(layer_0[1148] | layer_0[888]); 
    assign out[935] = layer_0[156]; 
    assign out[936] = ~(layer_0[814] ^ layer_0[296]); 
    assign out[937] = ~layer_0[1070]; 
    assign out[938] = ~layer_0[315]; 
    assign out[939] = layer_0[13] | layer_0[606]; 
    assign out[940] = layer_0[155]; 
    assign out[941] = ~layer_0[1272]; 
    assign out[942] = ~layer_0[804] | (layer_0[510] & layer_0[804]); 
    assign out[943] = ~layer_0[252]; 
    assign out[944] = layer_0[782]; 
    assign out[945] = layer_0[535]; 
    assign out[946] = ~layer_0[181]; 
    assign out[947] = ~layer_0[858] | (layer_0[1166] & layer_0[858]); 
    assign out[948] = layer_0[797]; 
    assign out[949] = ~layer_0[954] | (layer_0[954] & layer_0[279]); 
    assign out[950] = layer_0[1011] ^ layer_0[1153]; 
    assign out[951] = ~layer_0[938]; 
    assign out[952] = layer_0[1134] ^ layer_0[1047]; 
    assign out[953] = ~layer_0[520] | (layer_0[520] & layer_0[453]); 
    assign out[954] = ~layer_0[909]; 
    assign out[955] = ~layer_0[1227] | (layer_0[796] & layer_0[1227]); 
    assign out[956] = layer_0[1180] & ~layer_0[700]; 
    assign out[957] = layer_0[120] ^ layer_0[202]; 
    assign out[958] = layer_0[486] | layer_0[576]; 
    assign out[959] = ~layer_0[114]; 
    assign out[960] = layer_0[529] ^ layer_0[586]; 
    assign out[961] = ~layer_0[47] | (layer_0[47] & layer_0[359]); 
    assign out[962] = layer_0[835]; 
    assign out[963] = layer_0[731] & ~layer_0[356]; 
    assign out[964] = ~layer_0[319]; 
    assign out[965] = ~layer_0[1068] | (layer_0[15] & layer_0[1068]); 
    assign out[966] = ~(layer_0[522] & layer_0[548]); 
    assign out[967] = layer_0[903] & ~layer_0[390]; 
    assign out[968] = layer_0[463] ^ layer_0[834]; 
    assign out[969] = ~(layer_0[740] ^ layer_0[460]); 
    assign out[970] = ~layer_0[1121] | (layer_0[281] & layer_0[1121]); 
    assign out[971] = layer_0[321]; 
    assign out[972] = ~layer_0[204]; 
    assign out[973] = layer_0[389] ^ layer_0[690]; 
    assign out[974] = ~(layer_0[680] ^ layer_0[704]); 
    assign out[975] = layer_0[374] & ~layer_0[129]; 
    assign out[976] = layer_0[1118]; 
    assign out[977] = ~(layer_0[815] ^ layer_0[752]); 
    assign out[978] = layer_0[988] & ~layer_0[1031]; 
    assign out[979] = layer_0[416] & layer_0[702]; 
    assign out[980] = layer_0[712]; 
    assign out[981] = ~(layer_0[53] ^ layer_0[422]); 
    assign out[982] = ~(layer_0[625] | layer_0[484]); 
    assign out[983] = layer_0[247] ^ layer_0[567]; 
    assign out[984] = layer_0[64] & layer_0[308]; 
    assign out[985] = ~(layer_0[288] & layer_0[1145]); 
    assign out[986] = ~layer_0[470] | (layer_0[470] & layer_0[29]); 
    assign out[987] = layer_0[161] ^ layer_0[825]; 
    assign out[988] = layer_0[1142]; 
    assign out[989] = layer_0[771] ^ layer_0[137]; 
    assign out[990] = layer_0[257] ^ layer_0[585]; 
    assign out[991] = ~layer_0[1046] | (layer_0[1046] & layer_0[413]); 
    assign out[992] = ~(layer_0[267] & layer_0[732]); 
    assign out[993] = ~layer_0[1146]; 
    assign out[994] = layer_0[632] | layer_0[426]; 
    assign out[995] = ~(layer_0[1080] ^ layer_0[888]); 
    assign out[996] = ~(layer_0[767] ^ layer_0[766]); 
    assign out[997] = ~(layer_0[646] | layer_0[292]); 
    assign out[998] = layer_0[1265] ^ layer_0[812]; 
    assign out[999] = ~(layer_0[1066] ^ layer_0[12]); 
    assign out[1000] = ~(layer_0[201] ^ layer_0[30]); 
    assign out[1001] = ~layer_0[772]; 
    assign out[1002] = ~(layer_0[730] ^ layer_0[21]); 
    assign out[1003] = layer_0[2]; 
    assign out[1004] = ~layer_0[892] | (layer_0[510] & layer_0[892]); 
    assign out[1005] = layer_0[1021]; 
    assign out[1006] = ~(layer_0[410] & layer_0[218]); 
    assign out[1007] = ~(layer_0[1213] | layer_0[57]); 
    assign out[1008] = layer_0[175] ^ layer_0[531]; 
    assign out[1009] = ~layer_0[451] | (layer_0[451] & layer_0[856]); 
    assign out[1010] = ~layer_0[197]; 
    assign out[1011] = layer_0[818]; 
    assign out[1012] = ~(layer_0[75] | layer_0[103]); 
    assign out[1013] = ~(layer_0[611] | layer_0[1074]); 
    assign out[1014] = layer_0[129] ^ layer_0[686]; 
    assign out[1015] = layer_0[539]; 
    assign out[1016] = layer_0[406] ^ layer_0[152]; 
    assign out[1017] = layer_0[784] & layer_0[1175]; 
    assign out[1018] = ~(layer_0[875] | layer_0[934]); 
    assign out[1019] = ~(layer_0[1155] | layer_0[628]); 
    assign out[1020] = layer_0[1181] ^ layer_0[427]; 
    assign out[1021] = layer_0[417] & layer_0[1001]; 
    assign out[1022] = layer_0[1167]; 
    assign out[1023] = layer_0[730] & layer_0[1014]; 
    assign out[1024] = ~layer_0[1194]; 
    assign out[1025] = ~layer_0[925]; 
    assign out[1026] = layer_0[255] ^ layer_0[714]; 
    assign out[1027] = layer_0[1265]; 
    assign out[1028] = layer_0[776] & ~layer_0[853]; 
    assign out[1029] = ~(layer_0[326] ^ layer_0[543]); 
    assign out[1030] = ~(layer_0[1112] & layer_0[1032]); 
    assign out[1031] = ~layer_0[857]; 
    assign out[1032] = ~layer_0[884]; 
    assign out[1033] = ~(layer_0[1097] & layer_0[1160]); 
    assign out[1034] = layer_0[1244] ^ layer_0[535]; 
    assign out[1035] = ~(layer_0[1043] | layer_0[428]); 
    assign out[1036] = layer_0[651]; 
    assign out[1037] = layer_0[617] ^ layer_0[100]; 
    assign out[1038] = ~layer_0[868] | (layer_0[894] & layer_0[868]); 
    assign out[1039] = ~(layer_0[37] ^ layer_0[158]); 
    assign out[1040] = layer_0[38] & ~layer_0[857]; 
    assign out[1041] = ~(layer_0[179] | layer_0[169]); 
    assign out[1042] = layer_0[95]; 
    assign out[1043] = ~(layer_0[1043] | layer_0[196]); 
    assign out[1044] = layer_0[819] & ~layer_0[926]; 
    assign out[1045] = ~layer_0[1172]; 
    assign out[1046] = layer_0[922] | layer_0[59]; 
    assign out[1047] = layer_0[1254] | layer_0[1189]; 
    assign out[1048] = layer_0[217] & ~layer_0[1213]; 
    assign out[1049] = layer_0[1249]; 
    assign out[1050] = layer_0[1099]; 
    assign out[1051] = ~layer_0[991]; 
    assign out[1052] = layer_0[1149] | layer_0[461]; 
    assign out[1053] = layer_0[855] ^ layer_0[768]; 
    assign out[1054] = layer_0[1178]; 
    assign out[1055] = ~(layer_0[921] | layer_0[874]); 
    assign out[1056] = layer_0[589] & layer_0[383]; 
    assign out[1057] = ~(layer_0[832] ^ layer_0[977]); 
    assign out[1058] = layer_0[1125]; 
    assign out[1059] = ~layer_0[963]; 
    assign out[1060] = ~(layer_0[86] ^ layer_0[167]); 
    assign out[1061] = layer_0[854]; 
    assign out[1062] = layer_0[1180]; 
    assign out[1063] = layer_0[549] & layer_0[1264]; 
    assign out[1064] = layer_0[378] ^ layer_0[1133]; 
    assign out[1065] = layer_0[1035] ^ layer_0[499]; 
    assign out[1066] = ~layer_0[452]; 
    assign out[1067] = ~(layer_0[110] ^ layer_0[1266]); 
    assign out[1068] = ~layer_0[775]; 
    assign out[1069] = layer_0[532] & layer_0[408]; 
    assign out[1070] = layer_0[187] & layer_0[221]; 
    assign out[1071] = ~layer_0[612] | (layer_0[623] & layer_0[612]); 
    assign out[1072] = layer_0[634] ^ layer_0[421]; 
    assign out[1073] = layer_0[1041] ^ layer_0[420]; 
    assign out[1074] = ~(layer_0[980] ^ layer_0[543]); 
    assign out[1075] = ~(layer_0[431] ^ layer_0[377]); 
    assign out[1076] = layer_0[183] & ~layer_0[380]; 
    assign out[1077] = ~layer_0[845]; 
    assign out[1078] = layer_0[384] ^ layer_0[1060]; 
    assign out[1079] = layer_0[86] & ~layer_0[205]; 
    assign out[1080] = ~layer_0[1260] | (layer_0[210] & layer_0[1260]); 
    assign out[1081] = layer_0[272] & ~layer_0[921]; 
    assign out[1082] = layer_0[813] ^ layer_0[1236]; 
    assign out[1083] = layer_0[228] ^ layer_0[193]; 
    assign out[1084] = layer_0[870] & layer_0[50]; 
    assign out[1085] = layer_0[1279]; 
    assign out[1086] = layer_0[895]; 
    assign out[1087] = ~layer_0[837]; 
    assign out[1088] = ~(layer_0[639] ^ layer_0[211]); 
    assign out[1089] = ~(layer_0[881] ^ layer_0[852]); 
    assign out[1090] = ~layer_0[538]; 
    assign out[1091] = layer_0[401] & layer_0[396]; 
    assign out[1092] = layer_0[794] ^ layer_0[1239]; 
    assign out[1093] = layer_0[338]; 
    assign out[1094] = ~layer_0[1092] | (layer_0[1051] & layer_0[1092]); 
    assign out[1095] = layer_0[1171] ^ layer_0[94]; 
    assign out[1096] = layer_0[363] ^ layer_0[860]; 
    assign out[1097] = ~(layer_0[893] ^ layer_0[346]); 
    assign out[1098] = ~layer_0[760] | (layer_0[760] & layer_0[867]); 
    assign out[1099] = layer_0[233]; 
    assign out[1100] = ~(layer_0[399] & layer_0[1250]); 
    assign out[1101] = ~layer_0[830] | (layer_0[547] & layer_0[830]); 
    assign out[1102] = layer_0[474] ^ layer_0[759]; 
    assign out[1103] = ~(layer_0[354] | layer_0[322]); 
    assign out[1104] = ~(layer_0[231] ^ layer_0[1174]); 
    assign out[1105] = layer_0[1252] & ~layer_0[953]; 
    assign out[1106] = layer_0[652] & ~layer_0[300]; 
    assign out[1107] = ~(layer_0[542] | layer_0[800]); 
    assign out[1108] = layer_0[588] ^ layer_0[1102]; 
    assign out[1109] = layer_0[140] & layer_0[568]; 
    assign out[1110] = layer_0[363] & ~layer_0[484]; 
    assign out[1111] = layer_0[1096]; 
    assign out[1112] = ~layer_0[5]; 
    assign out[1113] = ~layer_0[479]; 
    assign out[1114] = layer_0[1152]; 
    assign out[1115] = ~(layer_0[809] ^ layer_0[163]); 
    assign out[1116] = layer_0[947] ^ layer_0[1042]; 
    assign out[1117] = layer_0[118] & ~layer_0[703]; 
    assign out[1118] = layer_0[1218] ^ layer_0[701]; 
    assign out[1119] = ~layer_0[125] | (layer_0[125] & layer_0[738]); 
    assign out[1120] = ~layer_0[1260]; 
    assign out[1121] = ~(layer_0[127] | layer_0[618]); 
    assign out[1122] = layer_0[1054] ^ layer_0[519]; 
    assign out[1123] = layer_0[593] & layer_0[9]; 
    assign out[1124] = layer_0[747] | layer_0[1234]; 
    assign out[1125] = layer_0[263]; 
    assign out[1126] = ~(layer_0[32] ^ layer_0[758]); 
    assign out[1127] = layer_0[511] ^ layer_0[766]; 
    assign out[1128] = layer_0[1064]; 
    assign out[1129] = layer_0[736]; 
    assign out[1130] = ~(layer_0[1113] ^ layer_0[553]); 
    assign out[1131] = ~(layer_0[228] ^ layer_0[336]); 
    assign out[1132] = layer_0[19] & layer_0[1026]; 
    assign out[1133] = ~layer_0[381] | (layer_0[541] & layer_0[381]); 
    assign out[1134] = ~(layer_0[1039] ^ layer_0[644]); 
    assign out[1135] = layer_0[1045] & ~layer_0[1215]; 
    assign out[1136] = ~layer_0[548] | (layer_0[548] & layer_0[799]); 
    assign out[1137] = ~(layer_0[1114] ^ layer_0[944]); 
    assign out[1138] = layer_0[77]; 
    assign out[1139] = layer_0[952] & ~layer_0[336]; 
    assign out[1140] = ~(layer_0[421] & layer_0[1205]); 
    assign out[1141] = layer_0[1128]; 
    assign out[1142] = ~layer_0[40] | (layer_0[40] & layer_0[545]); 
    assign out[1143] = ~layer_0[756]; 
    assign out[1144] = layer_0[581] ^ layer_0[1016]; 
    assign out[1145] = layer_0[495] & layer_0[578]; 
    assign out[1146] = layer_0[576] & ~layer_0[817]; 
    assign out[1147] = ~(layer_0[1005] ^ layer_0[782]); 
    assign out[1148] = layer_0[1218] & ~layer_0[1029]; 
    assign out[1149] = ~(layer_0[1267] ^ layer_0[502]); 
    assign out[1150] = ~(layer_0[933] | layer_0[772]); 
    assign out[1151] = layer_0[776] ^ layer_0[1228]; 
    assign out[1152] = ~layer_0[823]; 
    assign out[1153] = ~(layer_0[570] | layer_0[964]); 
    assign out[1154] = layer_0[815]; 
    assign out[1155] = layer_0[196] & ~layer_0[240]; 
    assign out[1156] = ~layer_0[97]; 
    assign out[1157] = layer_0[846] & ~layer_0[814]; 
    assign out[1158] = ~layer_0[655]; 
    assign out[1159] = ~layer_0[25]; 
    assign out[1160] = ~layer_0[529]; 
    assign out[1161] = layer_0[919] ^ layer_0[258]; 
    assign out[1162] = ~(layer_0[1035] ^ layer_0[833]); 
    assign out[1163] = ~(layer_0[876] ^ layer_0[1147]); 
    assign out[1164] = layer_0[956]; 
    assign out[1165] = layer_0[985] ^ layer_0[1130]; 
    assign out[1166] = layer_0[309]; 
    assign out[1167] = layer_0[764] | layer_0[996]; 
    assign out[1168] = layer_0[667] & ~layer_0[1177]; 
    assign out[1169] = layer_0[390] & layer_0[1012]; 
    assign out[1170] = ~layer_0[114]; 
    assign out[1171] = layer_0[391] & ~layer_0[176]; 
    assign out[1172] = ~(layer_0[905] ^ layer_0[154]); 
    assign out[1173] = layer_0[428]; 
    assign out[1174] = layer_0[997] & ~layer_0[51]; 
    assign out[1175] = layer_0[1256] & ~layer_0[910]; 
    assign out[1176] = layer_0[386] & layer_0[694]; 
    assign out[1177] = layer_0[540] & layer_0[1079]; 
    assign out[1178] = ~layer_0[785]; 
    assign out[1179] = layer_0[34] & ~layer_0[268]; 
    assign out[1180] = ~(layer_0[981] ^ layer_0[1040]); 
    assign out[1181] = layer_0[1111] & layer_0[1168]; 
    assign out[1182] = layer_0[454] & ~layer_0[262]; 
    assign out[1183] = ~layer_0[826]; 
    assign out[1184] = layer_0[901] ^ layer_0[162]; 
    assign out[1185] = ~layer_0[388]; 
    assign out[1186] = ~(layer_0[436] ^ layer_0[407]); 
    assign out[1187] = layer_0[991] & layer_0[1237]; 
    assign out[1188] = ~layer_0[61]; 
    assign out[1189] = ~(layer_0[120] & layer_0[481]); 
    assign out[1190] = layer_0[404] & ~layer_0[1228]; 
    assign out[1191] = layer_0[953] & layer_0[786]; 
    assign out[1192] = layer_0[331]; 
    assign out[1193] = ~layer_0[942]; 
    assign out[1194] = layer_0[99]; 
    assign out[1195] = layer_0[93] & ~layer_0[896]; 
    assign out[1196] = layer_0[708]; 
    assign out[1197] = layer_0[631] & ~layer_0[621]; 
    assign out[1198] = ~(layer_0[689] ^ layer_0[1146]); 
    assign out[1199] = ~(layer_0[1252] ^ layer_0[837]); 
    assign out[1200] = layer_0[665] & ~layer_0[459]; 
    assign out[1201] = layer_0[236]; 
    assign out[1202] = ~(layer_0[1106] ^ layer_0[689]); 
    assign out[1203] = layer_0[1045] & ~layer_0[574]; 
    assign out[1204] = ~(layer_0[791] ^ layer_0[193]); 
    assign out[1205] = ~layer_0[214]; 
    assign out[1206] = ~layer_0[83]; 
    assign out[1207] = layer_0[1258] & ~layer_0[697]; 
    assign out[1208] = ~(layer_0[505] & layer_0[483]); 
    assign out[1209] = layer_0[981]; 
    assign out[1210] = ~layer_0[232]; 
    assign out[1211] = layer_0[957]; 
    assign out[1212] = layer_0[691] ^ layer_0[450]; 
    assign out[1213] = layer_0[1270]; 
    assign out[1214] = layer_0[188] ^ layer_0[280]; 
    assign out[1215] = layer_0[990] & layer_0[728]; 
    assign out[1216] = layer_0[1236] ^ layer_0[828]; 
    assign out[1217] = ~layer_0[437] | (layer_0[73] & layer_0[437]); 
    assign out[1218] = layer_0[840] ^ layer_0[527]; 
    assign out[1219] = ~(layer_0[742] | layer_0[388]); 
    assign out[1220] = ~layer_0[302] | (layer_0[530] & layer_0[302]); 
    assign out[1221] = layer_0[884] ^ layer_0[1274]; 
    assign out[1222] = ~(layer_0[920] ^ layer_0[110]); 
    assign out[1223] = ~(layer_0[286] | layer_0[927]); 
    assign out[1224] = ~(layer_0[968] ^ layer_0[259]); 
    assign out[1225] = ~(layer_0[932] | layer_0[373]); 
    assign out[1226] = layer_0[69] ^ layer_0[1087]; 
    assign out[1227] = layer_0[1216] & layer_0[488]; 
    assign out[1228] = ~layer_0[961]; 
    assign out[1229] = ~layer_0[940]; 
    assign out[1230] = layer_0[995] & ~layer_0[1253]; 
    assign out[1231] = ~layer_0[1104] | (layer_0[1104] & layer_0[562]); 
    assign out[1232] = layer_0[536] & ~layer_0[713]; 
    assign out[1233] = layer_0[212] | layer_0[1012]; 
    assign out[1234] = layer_0[394] ^ layer_0[191]; 
    assign out[1235] = ~(layer_0[525] ^ layer_0[1173]); 
    assign out[1236] = layer_0[119]; 
    assign out[1237] = ~layer_0[166]; 
    assign out[1238] = ~(layer_0[1243] | layer_0[1181]); 
    assign out[1239] = layer_0[195] & ~layer_0[910]; 
    assign out[1240] = ~layer_0[1081] | (layer_0[875] & layer_0[1081]); 
    assign out[1241] = layer_0[236] & ~layer_0[993]; 
    assign out[1242] = layer_0[1088] & ~layer_0[803]; 
    assign out[1243] = layer_0[1038] & ~layer_0[771]; 
    assign out[1244] = layer_0[1072] ^ layer_0[1230]; 
    assign out[1245] = layer_0[1270] & ~layer_0[1039]; 
    assign out[1246] = layer_0[793]; 
    assign out[1247] = layer_0[908] & layer_0[971]; 
    assign out[1248] = ~(layer_0[158] ^ layer_0[96]); 
    assign out[1249] = ~(layer_0[262] & layer_0[653]); 
    assign out[1250] = ~layer_0[385]; 
    assign out[1251] = layer_0[426] & layer_0[902]; 
    assign out[1252] = ~(layer_0[72] ^ layer_0[316]); 
    assign out[1253] = ~(layer_0[1206] ^ layer_0[652]); 
    assign out[1254] = ~layer_0[319]; 
    assign out[1255] = ~(layer_0[49] ^ layer_0[741]); 
    assign out[1256] = layer_0[28] ^ layer_0[128]; 
    assign out[1257] = layer_0[1149] & ~layer_0[7]; 
    assign out[1258] = layer_0[224]; 
    assign out[1259] = layer_0[1008] & ~layer_0[290]; 
    assign out[1260] = layer_0[670] ^ layer_0[925]; 
    assign out[1261] = ~(layer_0[1277] ^ layer_0[948]); 
    assign out[1262] = ~layer_0[1186] | (layer_0[1186] & layer_0[816]); 
    assign out[1263] = ~(layer_0[589] | layer_0[1024]); 
    assign out[1264] = ~(layer_0[34] ^ layer_0[870]); 
    assign out[1265] = ~(layer_0[635] | layer_0[1132]); 
    assign out[1266] = layer_0[361] & ~layer_0[832]; 
    assign out[1267] = ~layer_0[1169]; 
    assign out[1268] = ~(layer_0[539] | layer_0[1116]); 
    assign out[1269] = layer_0[509] & ~layer_0[451]; 
    assign out[1270] = 1'b0; 
    assign out[1271] = 1'b0; 
    assign out[1272] = 1'b0; 
    assign out[1273] = 1'b0; 
    assign out[1274] = 1'b0; 
    assign out[1275] = 1'b0; 
    assign out[1276] = 1'b0; 
    assign out[1277] = 1'b0; 
    assign out[1278] = 1'b0; 
    assign out[1279] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[126:0] = out[126:0];
    assign categories[253:127] = out[254:128];
    assign categories[380:254] = out[382:256];
    assign categories[507:381] = out[510:384];
    assign categories[634:508] = out[638:512];
    assign categories[761:635] = out[766:640];
    assign categories[888:762] = out[894:768];
    assign categories[1015:889] = out[1022:896];
    assign categories[1142:1016] = out[1150:1024];
    assign categories[1269:1143] = out[1278:1152];

endmodule
