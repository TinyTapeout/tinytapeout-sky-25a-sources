magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -125 272 -67 278
rect 67 272 125 278
rect -125 238 -113 272
rect 67 238 79 272
rect -125 232 -67 238
rect 67 232 125 238
rect -221 -238 -163 -232
rect -29 -238 29 -232
rect 163 -238 221 -232
rect -221 -272 -209 -238
rect -29 -272 -17 -238
rect 163 -272 175 -238
rect -221 -278 -163 -272
rect -29 -278 29 -272
rect 163 -278 221 -272
<< pwell >>
rect -397 -400 397 400
<< nmos >>
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
<< ndiff >>
rect -269 187 -207 200
rect -269 153 -257 187
rect -223 153 -207 187
rect -269 119 -207 153
rect -269 85 -257 119
rect -223 85 -207 119
rect -269 51 -207 85
rect -269 17 -257 51
rect -223 17 -207 51
rect -269 -17 -207 17
rect -269 -51 -257 -17
rect -223 -51 -207 -17
rect -269 -85 -207 -51
rect -269 -119 -257 -85
rect -223 -119 -207 -85
rect -269 -153 -207 -119
rect -269 -187 -257 -153
rect -223 -187 -207 -153
rect -269 -200 -207 -187
rect -177 187 -111 200
rect -177 153 -161 187
rect -127 153 -111 187
rect -177 119 -111 153
rect -177 85 -161 119
rect -127 85 -111 119
rect -177 51 -111 85
rect -177 17 -161 51
rect -127 17 -111 51
rect -177 -17 -111 17
rect -177 -51 -161 -17
rect -127 -51 -111 -17
rect -177 -85 -111 -51
rect -177 -119 -161 -85
rect -127 -119 -111 -85
rect -177 -153 -111 -119
rect -177 -187 -161 -153
rect -127 -187 -111 -153
rect -177 -200 -111 -187
rect -81 187 -15 200
rect -81 153 -65 187
rect -31 153 -15 187
rect -81 119 -15 153
rect -81 85 -65 119
rect -31 85 -15 119
rect -81 51 -15 85
rect -81 17 -65 51
rect -31 17 -15 51
rect -81 -17 -15 17
rect -81 -51 -65 -17
rect -31 -51 -15 -17
rect -81 -85 -15 -51
rect -81 -119 -65 -85
rect -31 -119 -15 -85
rect -81 -153 -15 -119
rect -81 -187 -65 -153
rect -31 -187 -15 -153
rect -81 -200 -15 -187
rect 15 187 81 200
rect 15 153 31 187
rect 65 153 81 187
rect 15 119 81 153
rect 15 85 31 119
rect 65 85 81 119
rect 15 51 81 85
rect 15 17 31 51
rect 65 17 81 51
rect 15 -17 81 17
rect 15 -51 31 -17
rect 65 -51 81 -17
rect 15 -85 81 -51
rect 15 -119 31 -85
rect 65 -119 81 -85
rect 15 -153 81 -119
rect 15 -187 31 -153
rect 65 -187 81 -153
rect 15 -200 81 -187
rect 111 187 177 200
rect 111 153 127 187
rect 161 153 177 187
rect 111 119 177 153
rect 111 85 127 119
rect 161 85 177 119
rect 111 51 177 85
rect 111 17 127 51
rect 161 17 177 51
rect 111 -17 177 17
rect 111 -51 127 -17
rect 161 -51 177 -17
rect 111 -85 177 -51
rect 111 -119 127 -85
rect 161 -119 177 -85
rect 111 -153 177 -119
rect 111 -187 127 -153
rect 161 -187 177 -153
rect 111 -200 177 -187
rect 207 187 269 200
rect 207 153 223 187
rect 257 153 269 187
rect 207 119 269 153
rect 207 85 223 119
rect 257 85 269 119
rect 207 51 269 85
rect 207 17 223 51
rect 257 17 269 51
rect 207 -17 269 17
rect 207 -51 223 -17
rect 257 -51 269 -17
rect 207 -85 269 -51
rect 207 -119 223 -85
rect 257 -119 269 -85
rect 207 -153 269 -119
rect 207 -187 223 -153
rect 257 -187 269 -153
rect 207 -200 269 -187
<< ndiffc >>
rect -257 153 -223 187
rect -257 85 -223 119
rect -257 17 -223 51
rect -257 -51 -223 -17
rect -257 -119 -223 -85
rect -257 -187 -223 -153
rect -161 153 -127 187
rect -161 85 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -85
rect -161 -187 -127 -153
rect -65 153 -31 187
rect -65 85 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -85
rect -65 -187 -31 -153
rect 31 153 65 187
rect 31 85 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -85
rect 31 -187 65 -153
rect 127 153 161 187
rect 127 85 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -85
rect 127 -187 161 -153
rect 223 153 257 187
rect 223 85 257 119
rect 223 17 257 51
rect 223 -51 257 -17
rect 223 -119 257 -85
rect 223 -187 257 -153
<< psubdiff >>
rect -371 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 371 374
rect -371 255 -337 340
rect -371 187 -337 221
rect 337 255 371 340
rect -371 119 -337 153
rect -371 51 -337 85
rect -371 -17 -337 17
rect -371 -85 -337 -51
rect -371 -153 -337 -119
rect -371 -221 -337 -187
rect 337 187 371 221
rect 337 119 371 153
rect 337 51 371 85
rect 337 -17 371 17
rect 337 -85 371 -51
rect 337 -153 371 -119
rect -371 -340 -337 -255
rect 337 -221 371 -187
rect 337 -340 371 -255
rect -371 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 371 -340
<< psubdiffcont >>
rect -255 340 -221 374
rect -187 340 -153 374
rect -119 340 -85 374
rect -51 340 -17 374
rect 17 340 51 374
rect 85 340 119 374
rect 153 340 187 374
rect 221 340 255 374
rect -371 221 -337 255
rect 337 221 371 255
rect -371 153 -337 187
rect -371 85 -337 119
rect -371 17 -337 51
rect -371 -51 -337 -17
rect -371 -119 -337 -85
rect -371 -187 -337 -153
rect 337 153 371 187
rect 337 85 371 119
rect 337 17 371 51
rect 337 -51 371 -17
rect 337 -119 371 -85
rect 337 -187 371 -153
rect -371 -255 -337 -221
rect 337 -255 371 -221
rect -255 -374 -221 -340
rect -187 -374 -153 -340
rect -119 -374 -85 -340
rect -51 -374 -17 -340
rect 17 -374 51 -340
rect 85 -374 119 -340
rect 153 -374 187 -340
rect 221 -374 255 -340
<< poly >>
rect -129 272 -63 288
rect -129 238 -113 272
rect -79 238 -63 272
rect -207 200 -177 226
rect -129 222 -63 238
rect 63 272 129 288
rect 63 238 79 272
rect 113 238 129 272
rect -111 200 -81 222
rect -15 200 15 226
rect 63 222 129 238
rect 81 200 111 222
rect 177 200 207 226
rect -207 -222 -177 -200
rect -225 -238 -159 -222
rect -111 -226 -81 -200
rect -15 -222 15 -200
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -225 -288 -159 -272
rect -33 -238 33 -222
rect 81 -226 111 -200
rect 177 -222 207 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 159 -238 225 -222
rect 159 -272 175 -238
rect 209 -272 225 -238
rect 159 -288 225 -272
<< polycont >>
rect -113 238 -79 272
rect 79 238 113 272
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
<< locali >>
rect -371 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 371 374
rect -371 255 -337 340
rect -129 238 -113 272
rect -79 238 -63 272
rect 63 238 79 272
rect 113 238 129 272
rect 337 255 371 340
rect -371 187 -337 221
rect -371 119 -337 153
rect -371 51 -337 85
rect -371 -17 -337 17
rect -371 -85 -337 -51
rect -371 -153 -337 -119
rect -371 -221 -337 -187
rect -257 187 -223 204
rect -257 119 -223 127
rect -257 51 -223 55
rect -257 -55 -223 -51
rect -257 -127 -223 -119
rect -257 -204 -223 -187
rect -161 187 -127 204
rect -161 119 -127 127
rect -161 51 -127 55
rect -161 -55 -127 -51
rect -161 -127 -127 -119
rect -161 -204 -127 -187
rect -65 187 -31 204
rect -65 119 -31 127
rect -65 51 -31 55
rect -65 -55 -31 -51
rect -65 -127 -31 -119
rect -65 -204 -31 -187
rect 31 187 65 204
rect 31 119 65 127
rect 31 51 65 55
rect 31 -55 65 -51
rect 31 -127 65 -119
rect 31 -204 65 -187
rect 127 187 161 204
rect 127 119 161 127
rect 127 51 161 55
rect 127 -55 161 -51
rect 127 -127 161 -119
rect 127 -204 161 -187
rect 223 187 257 204
rect 223 119 257 127
rect 223 51 257 55
rect 223 -55 257 -51
rect 223 -127 257 -119
rect 223 -204 257 -187
rect 337 187 371 221
rect 337 119 371 153
rect 337 51 371 85
rect 337 -17 371 17
rect 337 -85 371 -51
rect 337 -153 371 -119
rect 337 -221 371 -187
rect -371 -340 -337 -255
rect -225 -272 -209 -238
rect -175 -272 -159 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 159 -272 175 -238
rect 209 -272 225 -238
rect 337 -340 371 -255
rect -371 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 371 -340
<< viali >>
rect -113 238 -79 272
rect 79 238 113 272
rect -257 153 -223 161
rect -257 127 -223 153
rect -257 85 -223 89
rect -257 55 -223 85
rect -257 -17 -223 17
rect -257 -85 -223 -55
rect -257 -89 -223 -85
rect -257 -153 -223 -127
rect -257 -161 -223 -153
rect -161 153 -127 161
rect -161 127 -127 153
rect -161 85 -127 89
rect -161 55 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -55
rect -161 -89 -127 -85
rect -161 -153 -127 -127
rect -161 -161 -127 -153
rect -65 153 -31 161
rect -65 127 -31 153
rect -65 85 -31 89
rect -65 55 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -55
rect -65 -89 -31 -85
rect -65 -153 -31 -127
rect -65 -161 -31 -153
rect 31 153 65 161
rect 31 127 65 153
rect 31 85 65 89
rect 31 55 65 85
rect 31 -17 65 17
rect 31 -85 65 -55
rect 31 -89 65 -85
rect 31 -153 65 -127
rect 31 -161 65 -153
rect 127 153 161 161
rect 127 127 161 153
rect 127 85 161 89
rect 127 55 161 85
rect 127 -17 161 17
rect 127 -85 161 -55
rect 127 -89 161 -85
rect 127 -153 161 -127
rect 127 -161 161 -153
rect 223 153 257 161
rect 223 127 257 153
rect 223 85 257 89
rect 223 55 257 85
rect 223 -17 257 17
rect 223 -85 257 -55
rect 223 -89 257 -85
rect 223 -153 257 -127
rect 223 -161 257 -153
rect -209 -272 -175 -238
rect -17 -272 17 -238
rect 175 -272 209 -238
<< metal1 >>
rect -125 272 -67 278
rect -125 238 -113 272
rect -79 238 -67 272
rect -125 232 -67 238
rect 67 272 125 278
rect 67 238 79 272
rect 113 238 125 272
rect 67 232 125 238
rect -263 161 -217 200
rect -263 127 -257 161
rect -223 127 -217 161
rect -263 89 -217 127
rect -263 55 -257 89
rect -223 55 -217 89
rect -263 17 -217 55
rect -263 -17 -257 17
rect -223 -17 -217 17
rect -263 -55 -217 -17
rect -263 -89 -257 -55
rect -223 -89 -217 -55
rect -263 -127 -217 -89
rect -263 -161 -257 -127
rect -223 -161 -217 -127
rect -263 -200 -217 -161
rect -167 161 -121 200
rect -167 127 -161 161
rect -127 127 -121 161
rect -167 89 -121 127
rect -167 55 -161 89
rect -127 55 -121 89
rect -167 17 -121 55
rect -167 -17 -161 17
rect -127 -17 -121 17
rect -167 -55 -121 -17
rect -167 -89 -161 -55
rect -127 -89 -121 -55
rect -167 -127 -121 -89
rect -167 -161 -161 -127
rect -127 -161 -121 -127
rect -167 -200 -121 -161
rect -71 161 -25 200
rect -71 127 -65 161
rect -31 127 -25 161
rect -71 89 -25 127
rect -71 55 -65 89
rect -31 55 -25 89
rect -71 17 -25 55
rect -71 -17 -65 17
rect -31 -17 -25 17
rect -71 -55 -25 -17
rect -71 -89 -65 -55
rect -31 -89 -25 -55
rect -71 -127 -25 -89
rect -71 -161 -65 -127
rect -31 -161 -25 -127
rect -71 -200 -25 -161
rect 25 161 71 200
rect 25 127 31 161
rect 65 127 71 161
rect 25 89 71 127
rect 25 55 31 89
rect 65 55 71 89
rect 25 17 71 55
rect 25 -17 31 17
rect 65 -17 71 17
rect 25 -55 71 -17
rect 25 -89 31 -55
rect 65 -89 71 -55
rect 25 -127 71 -89
rect 25 -161 31 -127
rect 65 -161 71 -127
rect 25 -200 71 -161
rect 121 161 167 200
rect 121 127 127 161
rect 161 127 167 161
rect 121 89 167 127
rect 121 55 127 89
rect 161 55 167 89
rect 121 17 167 55
rect 121 -17 127 17
rect 161 -17 167 17
rect 121 -55 167 -17
rect 121 -89 127 -55
rect 161 -89 167 -55
rect 121 -127 167 -89
rect 121 -161 127 -127
rect 161 -161 167 -127
rect 121 -200 167 -161
rect 217 161 263 200
rect 217 127 223 161
rect 257 127 263 161
rect 217 89 263 127
rect 217 55 223 89
rect 257 55 263 89
rect 217 17 263 55
rect 217 -17 223 17
rect 257 -17 263 17
rect 217 -55 263 -17
rect 217 -89 223 -55
rect 257 -89 263 -55
rect 217 -127 263 -89
rect 217 -161 223 -127
rect 257 -161 263 -127
rect 217 -200 263 -161
rect -221 -238 -163 -232
rect -221 -272 -209 -238
rect -175 -272 -163 -238
rect -221 -278 -163 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 163 -238 221 -232
rect 163 -272 175 -238
rect 209 -272 221 -238
rect 163 -278 221 -272
<< properties >>
string FIXED_BBOX -354 -357 354 357
<< end >>
