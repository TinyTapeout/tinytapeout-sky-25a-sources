magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -88 1572 -30 1578
rect 30 1572 88 1578
rect -88 1538 -76 1572
rect 30 1538 42 1572
rect -88 1532 -30 1538
rect 30 1532 88 1538
rect -88 -1538 -30 -1532
rect 30 -1538 88 -1532
rect -88 -1572 -76 -1538
rect 30 -1572 42 -1538
rect -88 -1578 -30 -1572
rect 30 -1578 88 -1572
<< pwell >>
rect -275 -1700 275 1700
<< nmos >>
rect -89 -1500 -29 1500
rect 29 -1500 89 1500
<< ndiff >>
rect -147 1479 -89 1500
rect -147 1445 -135 1479
rect -101 1445 -89 1479
rect -147 1411 -89 1445
rect -147 1377 -135 1411
rect -101 1377 -89 1411
rect -147 1343 -89 1377
rect -147 1309 -135 1343
rect -101 1309 -89 1343
rect -147 1275 -89 1309
rect -147 1241 -135 1275
rect -101 1241 -89 1275
rect -147 1207 -89 1241
rect -147 1173 -135 1207
rect -101 1173 -89 1207
rect -147 1139 -89 1173
rect -147 1105 -135 1139
rect -101 1105 -89 1139
rect -147 1071 -89 1105
rect -147 1037 -135 1071
rect -101 1037 -89 1071
rect -147 1003 -89 1037
rect -147 969 -135 1003
rect -101 969 -89 1003
rect -147 935 -89 969
rect -147 901 -135 935
rect -101 901 -89 935
rect -147 867 -89 901
rect -147 833 -135 867
rect -101 833 -89 867
rect -147 799 -89 833
rect -147 765 -135 799
rect -101 765 -89 799
rect -147 731 -89 765
rect -147 697 -135 731
rect -101 697 -89 731
rect -147 663 -89 697
rect -147 629 -135 663
rect -101 629 -89 663
rect -147 595 -89 629
rect -147 561 -135 595
rect -101 561 -89 595
rect -147 527 -89 561
rect -147 493 -135 527
rect -101 493 -89 527
rect -147 459 -89 493
rect -147 425 -135 459
rect -101 425 -89 459
rect -147 391 -89 425
rect -147 357 -135 391
rect -101 357 -89 391
rect -147 323 -89 357
rect -147 289 -135 323
rect -101 289 -89 323
rect -147 255 -89 289
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -289 -89 -255
rect -147 -323 -135 -289
rect -101 -323 -89 -289
rect -147 -357 -89 -323
rect -147 -391 -135 -357
rect -101 -391 -89 -357
rect -147 -425 -89 -391
rect -147 -459 -135 -425
rect -101 -459 -89 -425
rect -147 -493 -89 -459
rect -147 -527 -135 -493
rect -101 -527 -89 -493
rect -147 -561 -89 -527
rect -147 -595 -135 -561
rect -101 -595 -89 -561
rect -147 -629 -89 -595
rect -147 -663 -135 -629
rect -101 -663 -89 -629
rect -147 -697 -89 -663
rect -147 -731 -135 -697
rect -101 -731 -89 -697
rect -147 -765 -89 -731
rect -147 -799 -135 -765
rect -101 -799 -89 -765
rect -147 -833 -89 -799
rect -147 -867 -135 -833
rect -101 -867 -89 -833
rect -147 -901 -89 -867
rect -147 -935 -135 -901
rect -101 -935 -89 -901
rect -147 -969 -89 -935
rect -147 -1003 -135 -969
rect -101 -1003 -89 -969
rect -147 -1037 -89 -1003
rect -147 -1071 -135 -1037
rect -101 -1071 -89 -1037
rect -147 -1105 -89 -1071
rect -147 -1139 -135 -1105
rect -101 -1139 -89 -1105
rect -147 -1173 -89 -1139
rect -147 -1207 -135 -1173
rect -101 -1207 -89 -1173
rect -147 -1241 -89 -1207
rect -147 -1275 -135 -1241
rect -101 -1275 -89 -1241
rect -147 -1309 -89 -1275
rect -147 -1343 -135 -1309
rect -101 -1343 -89 -1309
rect -147 -1377 -89 -1343
rect -147 -1411 -135 -1377
rect -101 -1411 -89 -1377
rect -147 -1445 -89 -1411
rect -147 -1479 -135 -1445
rect -101 -1479 -89 -1445
rect -147 -1500 -89 -1479
rect -29 1479 29 1500
rect -29 1445 -17 1479
rect 17 1445 29 1479
rect -29 1411 29 1445
rect -29 1377 -17 1411
rect 17 1377 29 1411
rect -29 1343 29 1377
rect -29 1309 -17 1343
rect 17 1309 29 1343
rect -29 1275 29 1309
rect -29 1241 -17 1275
rect 17 1241 29 1275
rect -29 1207 29 1241
rect -29 1173 -17 1207
rect 17 1173 29 1207
rect -29 1139 29 1173
rect -29 1105 -17 1139
rect 17 1105 29 1139
rect -29 1071 29 1105
rect -29 1037 -17 1071
rect 17 1037 29 1071
rect -29 1003 29 1037
rect -29 969 -17 1003
rect 17 969 29 1003
rect -29 935 29 969
rect -29 901 -17 935
rect 17 901 29 935
rect -29 867 29 901
rect -29 833 -17 867
rect 17 833 29 867
rect -29 799 29 833
rect -29 765 -17 799
rect 17 765 29 799
rect -29 731 29 765
rect -29 697 -17 731
rect 17 697 29 731
rect -29 663 29 697
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -697 29 -663
rect -29 -731 -17 -697
rect 17 -731 29 -697
rect -29 -765 29 -731
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -833 29 -799
rect -29 -867 -17 -833
rect 17 -867 29 -833
rect -29 -901 29 -867
rect -29 -935 -17 -901
rect 17 -935 29 -901
rect -29 -969 29 -935
rect -29 -1003 -17 -969
rect 17 -1003 29 -969
rect -29 -1037 29 -1003
rect -29 -1071 -17 -1037
rect 17 -1071 29 -1037
rect -29 -1105 29 -1071
rect -29 -1139 -17 -1105
rect 17 -1139 29 -1105
rect -29 -1173 29 -1139
rect -29 -1207 -17 -1173
rect 17 -1207 29 -1173
rect -29 -1241 29 -1207
rect -29 -1275 -17 -1241
rect 17 -1275 29 -1241
rect -29 -1309 29 -1275
rect -29 -1343 -17 -1309
rect 17 -1343 29 -1309
rect -29 -1377 29 -1343
rect -29 -1411 -17 -1377
rect 17 -1411 29 -1377
rect -29 -1445 29 -1411
rect -29 -1479 -17 -1445
rect 17 -1479 29 -1445
rect -29 -1500 29 -1479
rect 89 1479 147 1500
rect 89 1445 101 1479
rect 135 1445 147 1479
rect 89 1411 147 1445
rect 89 1377 101 1411
rect 135 1377 147 1411
rect 89 1343 147 1377
rect 89 1309 101 1343
rect 135 1309 147 1343
rect 89 1275 147 1309
rect 89 1241 101 1275
rect 135 1241 147 1275
rect 89 1207 147 1241
rect 89 1173 101 1207
rect 135 1173 147 1207
rect 89 1139 147 1173
rect 89 1105 101 1139
rect 135 1105 147 1139
rect 89 1071 147 1105
rect 89 1037 101 1071
rect 135 1037 147 1071
rect 89 1003 147 1037
rect 89 969 101 1003
rect 135 969 147 1003
rect 89 935 147 969
rect 89 901 101 935
rect 135 901 147 935
rect 89 867 147 901
rect 89 833 101 867
rect 135 833 147 867
rect 89 799 147 833
rect 89 765 101 799
rect 135 765 147 799
rect 89 731 147 765
rect 89 697 101 731
rect 135 697 147 731
rect 89 663 147 697
rect 89 629 101 663
rect 135 629 147 663
rect 89 595 147 629
rect 89 561 101 595
rect 135 561 147 595
rect 89 527 147 561
rect 89 493 101 527
rect 135 493 147 527
rect 89 459 147 493
rect 89 425 101 459
rect 135 425 147 459
rect 89 391 147 425
rect 89 357 101 391
rect 135 357 147 391
rect 89 323 147 357
rect 89 289 101 323
rect 135 289 147 323
rect 89 255 147 289
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -289 147 -255
rect 89 -323 101 -289
rect 135 -323 147 -289
rect 89 -357 147 -323
rect 89 -391 101 -357
rect 135 -391 147 -357
rect 89 -425 147 -391
rect 89 -459 101 -425
rect 135 -459 147 -425
rect 89 -493 147 -459
rect 89 -527 101 -493
rect 135 -527 147 -493
rect 89 -561 147 -527
rect 89 -595 101 -561
rect 135 -595 147 -561
rect 89 -629 147 -595
rect 89 -663 101 -629
rect 135 -663 147 -629
rect 89 -697 147 -663
rect 89 -731 101 -697
rect 135 -731 147 -697
rect 89 -765 147 -731
rect 89 -799 101 -765
rect 135 -799 147 -765
rect 89 -833 147 -799
rect 89 -867 101 -833
rect 135 -867 147 -833
rect 89 -901 147 -867
rect 89 -935 101 -901
rect 135 -935 147 -901
rect 89 -969 147 -935
rect 89 -1003 101 -969
rect 135 -1003 147 -969
rect 89 -1037 147 -1003
rect 89 -1071 101 -1037
rect 135 -1071 147 -1037
rect 89 -1105 147 -1071
rect 89 -1139 101 -1105
rect 135 -1139 147 -1105
rect 89 -1173 147 -1139
rect 89 -1207 101 -1173
rect 135 -1207 147 -1173
rect 89 -1241 147 -1207
rect 89 -1275 101 -1241
rect 135 -1275 147 -1241
rect 89 -1309 147 -1275
rect 89 -1343 101 -1309
rect 135 -1343 147 -1309
rect 89 -1377 147 -1343
rect 89 -1411 101 -1377
rect 135 -1411 147 -1377
rect 89 -1445 147 -1411
rect 89 -1479 101 -1445
rect 135 -1479 147 -1445
rect 89 -1500 147 -1479
<< ndiffc >>
rect -135 1445 -101 1479
rect -135 1377 -101 1411
rect -135 1309 -101 1343
rect -135 1241 -101 1275
rect -135 1173 -101 1207
rect -135 1105 -101 1139
rect -135 1037 -101 1071
rect -135 969 -101 1003
rect -135 901 -101 935
rect -135 833 -101 867
rect -135 765 -101 799
rect -135 697 -101 731
rect -135 629 -101 663
rect -135 561 -101 595
rect -135 493 -101 527
rect -135 425 -101 459
rect -135 357 -101 391
rect -135 289 -101 323
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -135 -323 -101 -289
rect -135 -391 -101 -357
rect -135 -459 -101 -425
rect -135 -527 -101 -493
rect -135 -595 -101 -561
rect -135 -663 -101 -629
rect -135 -731 -101 -697
rect -135 -799 -101 -765
rect -135 -867 -101 -833
rect -135 -935 -101 -901
rect -135 -1003 -101 -969
rect -135 -1071 -101 -1037
rect -135 -1139 -101 -1105
rect -135 -1207 -101 -1173
rect -135 -1275 -101 -1241
rect -135 -1343 -101 -1309
rect -135 -1411 -101 -1377
rect -135 -1479 -101 -1445
rect -17 1445 17 1479
rect -17 1377 17 1411
rect -17 1309 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1139
rect -17 1037 17 1071
rect -17 969 17 1003
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1003 17 -969
rect -17 -1071 17 -1037
rect -17 -1139 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1309
rect -17 -1411 17 -1377
rect -17 -1479 17 -1445
rect 101 1445 135 1479
rect 101 1377 135 1411
rect 101 1309 135 1343
rect 101 1241 135 1275
rect 101 1173 135 1207
rect 101 1105 135 1139
rect 101 1037 135 1071
rect 101 969 135 1003
rect 101 901 135 935
rect 101 833 135 867
rect 101 765 135 799
rect 101 697 135 731
rect 101 629 135 663
rect 101 561 135 595
rect 101 493 135 527
rect 101 425 135 459
rect 101 357 135 391
rect 101 289 135 323
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
rect 101 -323 135 -289
rect 101 -391 135 -357
rect 101 -459 135 -425
rect 101 -527 135 -493
rect 101 -595 135 -561
rect 101 -663 135 -629
rect 101 -731 135 -697
rect 101 -799 135 -765
rect 101 -867 135 -833
rect 101 -935 135 -901
rect 101 -1003 135 -969
rect 101 -1071 135 -1037
rect 101 -1139 135 -1105
rect 101 -1207 135 -1173
rect 101 -1275 135 -1241
rect 101 -1343 135 -1309
rect 101 -1411 135 -1377
rect 101 -1479 135 -1445
<< psubdiff >>
rect -249 1640 -153 1674
rect -119 1640 -85 1674
rect -51 1640 -17 1674
rect 17 1640 51 1674
rect 85 1640 119 1674
rect 153 1640 249 1674
rect -249 1547 -215 1640
rect 215 1547 249 1640
rect -249 1479 -215 1513
rect -249 1411 -215 1445
rect -249 1343 -215 1377
rect -249 1275 -215 1309
rect -249 1207 -215 1241
rect -249 1139 -215 1173
rect -249 1071 -215 1105
rect -249 1003 -215 1037
rect -249 935 -215 969
rect -249 867 -215 901
rect -249 799 -215 833
rect -249 731 -215 765
rect -249 663 -215 697
rect -249 595 -215 629
rect -249 527 -215 561
rect -249 459 -215 493
rect -249 391 -215 425
rect -249 323 -215 357
rect -249 255 -215 289
rect -249 187 -215 221
rect -249 119 -215 153
rect -249 51 -215 85
rect -249 -17 -215 17
rect -249 -85 -215 -51
rect -249 -153 -215 -119
rect -249 -221 -215 -187
rect -249 -289 -215 -255
rect -249 -357 -215 -323
rect -249 -425 -215 -391
rect -249 -493 -215 -459
rect -249 -561 -215 -527
rect -249 -629 -215 -595
rect -249 -697 -215 -663
rect -249 -765 -215 -731
rect -249 -833 -215 -799
rect -249 -901 -215 -867
rect -249 -969 -215 -935
rect -249 -1037 -215 -1003
rect -249 -1105 -215 -1071
rect -249 -1173 -215 -1139
rect -249 -1241 -215 -1207
rect -249 -1309 -215 -1275
rect -249 -1377 -215 -1343
rect -249 -1445 -215 -1411
rect -249 -1513 -215 -1479
rect 215 1479 249 1513
rect 215 1411 249 1445
rect 215 1343 249 1377
rect 215 1275 249 1309
rect 215 1207 249 1241
rect 215 1139 249 1173
rect 215 1071 249 1105
rect 215 1003 249 1037
rect 215 935 249 969
rect 215 867 249 901
rect 215 799 249 833
rect 215 731 249 765
rect 215 663 249 697
rect 215 595 249 629
rect 215 527 249 561
rect 215 459 249 493
rect 215 391 249 425
rect 215 323 249 357
rect 215 255 249 289
rect 215 187 249 221
rect 215 119 249 153
rect 215 51 249 85
rect 215 -17 249 17
rect 215 -85 249 -51
rect 215 -153 249 -119
rect 215 -221 249 -187
rect 215 -289 249 -255
rect 215 -357 249 -323
rect 215 -425 249 -391
rect 215 -493 249 -459
rect 215 -561 249 -527
rect 215 -629 249 -595
rect 215 -697 249 -663
rect 215 -765 249 -731
rect 215 -833 249 -799
rect 215 -901 249 -867
rect 215 -969 249 -935
rect 215 -1037 249 -1003
rect 215 -1105 249 -1071
rect 215 -1173 249 -1139
rect 215 -1241 249 -1207
rect 215 -1309 249 -1275
rect 215 -1377 249 -1343
rect 215 -1445 249 -1411
rect 215 -1513 249 -1479
rect -249 -1640 -215 -1547
rect 215 -1640 249 -1547
rect -249 -1674 -153 -1640
rect -119 -1674 -85 -1640
rect -51 -1674 -17 -1640
rect 17 -1674 51 -1640
rect 85 -1674 119 -1640
rect 153 -1674 249 -1640
<< psubdiffcont >>
rect -153 1640 -119 1674
rect -85 1640 -51 1674
rect -17 1640 17 1674
rect 51 1640 85 1674
rect 119 1640 153 1674
rect -249 1513 -215 1547
rect 215 1513 249 1547
rect -249 1445 -215 1479
rect -249 1377 -215 1411
rect -249 1309 -215 1343
rect -249 1241 -215 1275
rect -249 1173 -215 1207
rect -249 1105 -215 1139
rect -249 1037 -215 1071
rect -249 969 -215 1003
rect -249 901 -215 935
rect -249 833 -215 867
rect -249 765 -215 799
rect -249 697 -215 731
rect -249 629 -215 663
rect -249 561 -215 595
rect -249 493 -215 527
rect -249 425 -215 459
rect -249 357 -215 391
rect -249 289 -215 323
rect -249 221 -215 255
rect -249 153 -215 187
rect -249 85 -215 119
rect -249 17 -215 51
rect -249 -51 -215 -17
rect -249 -119 -215 -85
rect -249 -187 -215 -153
rect -249 -255 -215 -221
rect -249 -323 -215 -289
rect -249 -391 -215 -357
rect -249 -459 -215 -425
rect -249 -527 -215 -493
rect -249 -595 -215 -561
rect -249 -663 -215 -629
rect -249 -731 -215 -697
rect -249 -799 -215 -765
rect -249 -867 -215 -833
rect -249 -935 -215 -901
rect -249 -1003 -215 -969
rect -249 -1071 -215 -1037
rect -249 -1139 -215 -1105
rect -249 -1207 -215 -1173
rect -249 -1275 -215 -1241
rect -249 -1343 -215 -1309
rect -249 -1411 -215 -1377
rect -249 -1479 -215 -1445
rect 215 1445 249 1479
rect 215 1377 249 1411
rect 215 1309 249 1343
rect 215 1241 249 1275
rect 215 1173 249 1207
rect 215 1105 249 1139
rect 215 1037 249 1071
rect 215 969 249 1003
rect 215 901 249 935
rect 215 833 249 867
rect 215 765 249 799
rect 215 697 249 731
rect 215 629 249 663
rect 215 561 249 595
rect 215 493 249 527
rect 215 425 249 459
rect 215 357 249 391
rect 215 289 249 323
rect 215 221 249 255
rect 215 153 249 187
rect 215 85 249 119
rect 215 17 249 51
rect 215 -51 249 -17
rect 215 -119 249 -85
rect 215 -187 249 -153
rect 215 -255 249 -221
rect 215 -323 249 -289
rect 215 -391 249 -357
rect 215 -459 249 -425
rect 215 -527 249 -493
rect 215 -595 249 -561
rect 215 -663 249 -629
rect 215 -731 249 -697
rect 215 -799 249 -765
rect 215 -867 249 -833
rect 215 -935 249 -901
rect 215 -1003 249 -969
rect 215 -1071 249 -1037
rect 215 -1139 249 -1105
rect 215 -1207 249 -1173
rect 215 -1275 249 -1241
rect 215 -1343 249 -1309
rect 215 -1411 249 -1377
rect 215 -1479 249 -1445
rect -249 -1547 -215 -1513
rect 215 -1547 249 -1513
rect -153 -1674 -119 -1640
rect -85 -1674 -51 -1640
rect -17 -1674 17 -1640
rect 51 -1674 85 -1640
rect 119 -1674 153 -1640
<< poly >>
rect -92 1572 -26 1588
rect -92 1538 -76 1572
rect -42 1538 -26 1572
rect -92 1522 -26 1538
rect 26 1572 92 1588
rect 26 1538 42 1572
rect 76 1538 92 1572
rect 26 1522 92 1538
rect -89 1500 -29 1522
rect 29 1500 89 1522
rect -89 -1522 -29 -1500
rect 29 -1522 89 -1500
rect -92 -1538 -26 -1522
rect -92 -1572 -76 -1538
rect -42 -1572 -26 -1538
rect -92 -1588 -26 -1572
rect 26 -1538 92 -1522
rect 26 -1572 42 -1538
rect 76 -1572 92 -1538
rect 26 -1588 92 -1572
<< polycont >>
rect -76 1538 -42 1572
rect 42 1538 76 1572
rect -76 -1572 -42 -1538
rect 42 -1572 76 -1538
<< locali >>
rect -249 1640 -153 1674
rect -119 1640 -85 1674
rect -51 1640 -17 1674
rect 17 1640 51 1674
rect 85 1640 119 1674
rect 153 1640 249 1674
rect -249 1547 -215 1640
rect -92 1538 -76 1572
rect -42 1538 -26 1572
rect 26 1538 42 1572
rect 76 1538 92 1572
rect 215 1547 249 1640
rect -249 1479 -215 1513
rect -249 1411 -215 1445
rect -249 1343 -215 1377
rect -249 1275 -215 1309
rect -249 1207 -215 1241
rect -249 1139 -215 1173
rect -249 1071 -215 1105
rect -249 1003 -215 1037
rect -249 935 -215 969
rect -249 867 -215 901
rect -249 799 -215 833
rect -249 731 -215 765
rect -249 663 -215 697
rect -249 595 -215 629
rect -249 527 -215 561
rect -249 459 -215 493
rect -249 391 -215 425
rect -249 323 -215 357
rect -249 255 -215 289
rect -249 187 -215 221
rect -249 119 -215 153
rect -249 51 -215 85
rect -249 -17 -215 17
rect -249 -85 -215 -51
rect -249 -153 -215 -119
rect -249 -221 -215 -187
rect -249 -289 -215 -255
rect -249 -357 -215 -323
rect -249 -425 -215 -391
rect -249 -493 -215 -459
rect -249 -561 -215 -527
rect -249 -629 -215 -595
rect -249 -697 -215 -663
rect -249 -765 -215 -731
rect -249 -833 -215 -799
rect -249 -901 -215 -867
rect -249 -969 -215 -935
rect -249 -1037 -215 -1003
rect -249 -1105 -215 -1071
rect -249 -1173 -215 -1139
rect -249 -1241 -215 -1207
rect -249 -1309 -215 -1275
rect -249 -1377 -215 -1343
rect -249 -1445 -215 -1411
rect -249 -1513 -215 -1479
rect -135 1479 -101 1504
rect -135 1411 -101 1423
rect -135 1343 -101 1351
rect -135 1275 -101 1279
rect -135 1169 -101 1173
rect -135 1097 -101 1105
rect -135 1025 -101 1037
rect -135 953 -101 969
rect -135 881 -101 901
rect -135 809 -101 833
rect -135 737 -101 765
rect -135 665 -101 697
rect -135 595 -101 629
rect -135 527 -101 559
rect -135 459 -101 487
rect -135 391 -101 415
rect -135 323 -101 343
rect -135 255 -101 271
rect -135 187 -101 199
rect -135 119 -101 127
rect -135 51 -101 55
rect -135 -55 -101 -51
rect -135 -127 -101 -119
rect -135 -199 -101 -187
rect -135 -271 -101 -255
rect -135 -343 -101 -323
rect -135 -415 -101 -391
rect -135 -487 -101 -459
rect -135 -559 -101 -527
rect -135 -629 -101 -595
rect -135 -697 -101 -665
rect -135 -765 -101 -737
rect -135 -833 -101 -809
rect -135 -901 -101 -881
rect -135 -969 -101 -953
rect -135 -1037 -101 -1025
rect -135 -1105 -101 -1097
rect -135 -1173 -101 -1169
rect -135 -1279 -101 -1275
rect -135 -1351 -101 -1343
rect -135 -1423 -101 -1411
rect -135 -1504 -101 -1479
rect -17 1479 17 1504
rect -17 1411 17 1423
rect -17 1343 17 1351
rect -17 1275 17 1279
rect -17 1169 17 1173
rect -17 1097 17 1105
rect -17 1025 17 1037
rect -17 953 17 969
rect -17 881 17 901
rect -17 809 17 833
rect -17 737 17 765
rect -17 665 17 697
rect -17 595 17 629
rect -17 527 17 559
rect -17 459 17 487
rect -17 391 17 415
rect -17 323 17 343
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -343 17 -323
rect -17 -415 17 -391
rect -17 -487 17 -459
rect -17 -559 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -665
rect -17 -765 17 -737
rect -17 -833 17 -809
rect -17 -901 17 -881
rect -17 -969 17 -953
rect -17 -1037 17 -1025
rect -17 -1105 17 -1097
rect -17 -1173 17 -1169
rect -17 -1279 17 -1275
rect -17 -1351 17 -1343
rect -17 -1423 17 -1411
rect -17 -1504 17 -1479
rect 101 1479 135 1504
rect 101 1411 135 1423
rect 101 1343 135 1351
rect 101 1275 135 1279
rect 101 1169 135 1173
rect 101 1097 135 1105
rect 101 1025 135 1037
rect 101 953 135 969
rect 101 881 135 901
rect 101 809 135 833
rect 101 737 135 765
rect 101 665 135 697
rect 101 595 135 629
rect 101 527 135 559
rect 101 459 135 487
rect 101 391 135 415
rect 101 323 135 343
rect 101 255 135 271
rect 101 187 135 199
rect 101 119 135 127
rect 101 51 135 55
rect 101 -55 135 -51
rect 101 -127 135 -119
rect 101 -199 135 -187
rect 101 -271 135 -255
rect 101 -343 135 -323
rect 101 -415 135 -391
rect 101 -487 135 -459
rect 101 -559 135 -527
rect 101 -629 135 -595
rect 101 -697 135 -665
rect 101 -765 135 -737
rect 101 -833 135 -809
rect 101 -901 135 -881
rect 101 -969 135 -953
rect 101 -1037 135 -1025
rect 101 -1105 135 -1097
rect 101 -1173 135 -1169
rect 101 -1279 135 -1275
rect 101 -1351 135 -1343
rect 101 -1423 135 -1411
rect 101 -1504 135 -1479
rect 215 1479 249 1513
rect 215 1411 249 1445
rect 215 1343 249 1377
rect 215 1275 249 1309
rect 215 1207 249 1241
rect 215 1139 249 1173
rect 215 1071 249 1105
rect 215 1003 249 1037
rect 215 935 249 969
rect 215 867 249 901
rect 215 799 249 833
rect 215 731 249 765
rect 215 663 249 697
rect 215 595 249 629
rect 215 527 249 561
rect 215 459 249 493
rect 215 391 249 425
rect 215 323 249 357
rect 215 255 249 289
rect 215 187 249 221
rect 215 119 249 153
rect 215 51 249 85
rect 215 -17 249 17
rect 215 -85 249 -51
rect 215 -153 249 -119
rect 215 -221 249 -187
rect 215 -289 249 -255
rect 215 -357 249 -323
rect 215 -425 249 -391
rect 215 -493 249 -459
rect 215 -561 249 -527
rect 215 -629 249 -595
rect 215 -697 249 -663
rect 215 -765 249 -731
rect 215 -833 249 -799
rect 215 -901 249 -867
rect 215 -969 249 -935
rect 215 -1037 249 -1003
rect 215 -1105 249 -1071
rect 215 -1173 249 -1139
rect 215 -1241 249 -1207
rect 215 -1309 249 -1275
rect 215 -1377 249 -1343
rect 215 -1445 249 -1411
rect 215 -1513 249 -1479
rect -249 -1640 -215 -1547
rect -92 -1572 -76 -1538
rect -42 -1572 -26 -1538
rect 26 -1572 42 -1538
rect 76 -1572 92 -1538
rect 215 -1640 249 -1547
rect -249 -1674 -153 -1640
rect -119 -1674 -85 -1640
rect -51 -1674 -17 -1640
rect 17 -1674 51 -1640
rect 85 -1674 119 -1640
rect 153 -1674 249 -1640
<< viali >>
rect -76 1538 -42 1572
rect 42 1538 76 1572
rect -135 1445 -101 1457
rect -135 1423 -101 1445
rect -135 1377 -101 1385
rect -135 1351 -101 1377
rect -135 1309 -101 1313
rect -135 1279 -101 1309
rect -135 1207 -101 1241
rect -135 1139 -101 1169
rect -135 1135 -101 1139
rect -135 1071 -101 1097
rect -135 1063 -101 1071
rect -135 1003 -101 1025
rect -135 991 -101 1003
rect -135 935 -101 953
rect -135 919 -101 935
rect -135 867 -101 881
rect -135 847 -101 867
rect -135 799 -101 809
rect -135 775 -101 799
rect -135 731 -101 737
rect -135 703 -101 731
rect -135 663 -101 665
rect -135 631 -101 663
rect -135 561 -101 593
rect -135 559 -101 561
rect -135 493 -101 521
rect -135 487 -101 493
rect -135 425 -101 449
rect -135 415 -101 425
rect -135 357 -101 377
rect -135 343 -101 357
rect -135 289 -101 305
rect -135 271 -101 289
rect -135 221 -101 233
rect -135 199 -101 221
rect -135 153 -101 161
rect -135 127 -101 153
rect -135 85 -101 89
rect -135 55 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -55
rect -135 -89 -101 -85
rect -135 -153 -101 -127
rect -135 -161 -101 -153
rect -135 -221 -101 -199
rect -135 -233 -101 -221
rect -135 -289 -101 -271
rect -135 -305 -101 -289
rect -135 -357 -101 -343
rect -135 -377 -101 -357
rect -135 -425 -101 -415
rect -135 -449 -101 -425
rect -135 -493 -101 -487
rect -135 -521 -101 -493
rect -135 -561 -101 -559
rect -135 -593 -101 -561
rect -135 -663 -101 -631
rect -135 -665 -101 -663
rect -135 -731 -101 -703
rect -135 -737 -101 -731
rect -135 -799 -101 -775
rect -135 -809 -101 -799
rect -135 -867 -101 -847
rect -135 -881 -101 -867
rect -135 -935 -101 -919
rect -135 -953 -101 -935
rect -135 -1003 -101 -991
rect -135 -1025 -101 -1003
rect -135 -1071 -101 -1063
rect -135 -1097 -101 -1071
rect -135 -1139 -101 -1135
rect -135 -1169 -101 -1139
rect -135 -1241 -101 -1207
rect -135 -1309 -101 -1279
rect -135 -1313 -101 -1309
rect -135 -1377 -101 -1351
rect -135 -1385 -101 -1377
rect -135 -1445 -101 -1423
rect -135 -1457 -101 -1445
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect 101 1445 135 1457
rect 101 1423 135 1445
rect 101 1377 135 1385
rect 101 1351 135 1377
rect 101 1309 135 1313
rect 101 1279 135 1309
rect 101 1207 135 1241
rect 101 1139 135 1169
rect 101 1135 135 1139
rect 101 1071 135 1097
rect 101 1063 135 1071
rect 101 1003 135 1025
rect 101 991 135 1003
rect 101 935 135 953
rect 101 919 135 935
rect 101 867 135 881
rect 101 847 135 867
rect 101 799 135 809
rect 101 775 135 799
rect 101 731 135 737
rect 101 703 135 731
rect 101 663 135 665
rect 101 631 135 663
rect 101 561 135 593
rect 101 559 135 561
rect 101 493 135 521
rect 101 487 135 493
rect 101 425 135 449
rect 101 415 135 425
rect 101 357 135 377
rect 101 343 135 357
rect 101 289 135 305
rect 101 271 135 289
rect 101 221 135 233
rect 101 199 135 221
rect 101 153 135 161
rect 101 127 135 153
rect 101 85 135 89
rect 101 55 135 85
rect 101 -17 135 17
rect 101 -85 135 -55
rect 101 -89 135 -85
rect 101 -153 135 -127
rect 101 -161 135 -153
rect 101 -221 135 -199
rect 101 -233 135 -221
rect 101 -289 135 -271
rect 101 -305 135 -289
rect 101 -357 135 -343
rect 101 -377 135 -357
rect 101 -425 135 -415
rect 101 -449 135 -425
rect 101 -493 135 -487
rect 101 -521 135 -493
rect 101 -561 135 -559
rect 101 -593 135 -561
rect 101 -663 135 -631
rect 101 -665 135 -663
rect 101 -731 135 -703
rect 101 -737 135 -731
rect 101 -799 135 -775
rect 101 -809 135 -799
rect 101 -867 135 -847
rect 101 -881 135 -867
rect 101 -935 135 -919
rect 101 -953 135 -935
rect 101 -1003 135 -991
rect 101 -1025 135 -1003
rect 101 -1071 135 -1063
rect 101 -1097 135 -1071
rect 101 -1139 135 -1135
rect 101 -1169 135 -1139
rect 101 -1241 135 -1207
rect 101 -1309 135 -1279
rect 101 -1313 135 -1309
rect 101 -1377 135 -1351
rect 101 -1385 135 -1377
rect 101 -1445 135 -1423
rect 101 -1457 135 -1445
rect -76 -1572 -42 -1538
rect 42 -1572 76 -1538
<< metal1 >>
rect -88 1572 -30 1578
rect -88 1538 -76 1572
rect -42 1538 -30 1572
rect -88 1532 -30 1538
rect 30 1572 88 1578
rect 30 1538 42 1572
rect 76 1538 88 1572
rect 30 1532 88 1538
rect -141 1457 -95 1500
rect -141 1423 -135 1457
rect -101 1423 -95 1457
rect -141 1385 -95 1423
rect -141 1351 -135 1385
rect -101 1351 -95 1385
rect -141 1313 -95 1351
rect -141 1279 -135 1313
rect -101 1279 -95 1313
rect -141 1241 -95 1279
rect -141 1207 -135 1241
rect -101 1207 -95 1241
rect -141 1169 -95 1207
rect -141 1135 -135 1169
rect -101 1135 -95 1169
rect -141 1097 -95 1135
rect -141 1063 -135 1097
rect -101 1063 -95 1097
rect -141 1025 -95 1063
rect -141 991 -135 1025
rect -101 991 -95 1025
rect -141 953 -95 991
rect -141 919 -135 953
rect -101 919 -95 953
rect -141 881 -95 919
rect -141 847 -135 881
rect -101 847 -95 881
rect -141 809 -95 847
rect -141 775 -135 809
rect -101 775 -95 809
rect -141 737 -95 775
rect -141 703 -135 737
rect -101 703 -95 737
rect -141 665 -95 703
rect -141 631 -135 665
rect -101 631 -95 665
rect -141 593 -95 631
rect -141 559 -135 593
rect -101 559 -95 593
rect -141 521 -95 559
rect -141 487 -135 521
rect -101 487 -95 521
rect -141 449 -95 487
rect -141 415 -135 449
rect -101 415 -95 449
rect -141 377 -95 415
rect -141 343 -135 377
rect -101 343 -95 377
rect -141 305 -95 343
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -343 -95 -305
rect -141 -377 -135 -343
rect -101 -377 -95 -343
rect -141 -415 -95 -377
rect -141 -449 -135 -415
rect -101 -449 -95 -415
rect -141 -487 -95 -449
rect -141 -521 -135 -487
rect -101 -521 -95 -487
rect -141 -559 -95 -521
rect -141 -593 -135 -559
rect -101 -593 -95 -559
rect -141 -631 -95 -593
rect -141 -665 -135 -631
rect -101 -665 -95 -631
rect -141 -703 -95 -665
rect -141 -737 -135 -703
rect -101 -737 -95 -703
rect -141 -775 -95 -737
rect -141 -809 -135 -775
rect -101 -809 -95 -775
rect -141 -847 -95 -809
rect -141 -881 -135 -847
rect -101 -881 -95 -847
rect -141 -919 -95 -881
rect -141 -953 -135 -919
rect -101 -953 -95 -919
rect -141 -991 -95 -953
rect -141 -1025 -135 -991
rect -101 -1025 -95 -991
rect -141 -1063 -95 -1025
rect -141 -1097 -135 -1063
rect -101 -1097 -95 -1063
rect -141 -1135 -95 -1097
rect -141 -1169 -135 -1135
rect -101 -1169 -95 -1135
rect -141 -1207 -95 -1169
rect -141 -1241 -135 -1207
rect -101 -1241 -95 -1207
rect -141 -1279 -95 -1241
rect -141 -1313 -135 -1279
rect -101 -1313 -95 -1279
rect -141 -1351 -95 -1313
rect -141 -1385 -135 -1351
rect -101 -1385 -95 -1351
rect -141 -1423 -95 -1385
rect -141 -1457 -135 -1423
rect -101 -1457 -95 -1423
rect -141 -1500 -95 -1457
rect -23 1457 23 1500
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1500 23 -1457
rect 95 1457 141 1500
rect 95 1423 101 1457
rect 135 1423 141 1457
rect 95 1385 141 1423
rect 95 1351 101 1385
rect 135 1351 141 1385
rect 95 1313 141 1351
rect 95 1279 101 1313
rect 135 1279 141 1313
rect 95 1241 141 1279
rect 95 1207 101 1241
rect 135 1207 141 1241
rect 95 1169 141 1207
rect 95 1135 101 1169
rect 135 1135 141 1169
rect 95 1097 141 1135
rect 95 1063 101 1097
rect 135 1063 141 1097
rect 95 1025 141 1063
rect 95 991 101 1025
rect 135 991 141 1025
rect 95 953 141 991
rect 95 919 101 953
rect 135 919 141 953
rect 95 881 141 919
rect 95 847 101 881
rect 135 847 141 881
rect 95 809 141 847
rect 95 775 101 809
rect 135 775 141 809
rect 95 737 141 775
rect 95 703 101 737
rect 135 703 141 737
rect 95 665 141 703
rect 95 631 101 665
rect 135 631 141 665
rect 95 593 141 631
rect 95 559 101 593
rect 135 559 141 593
rect 95 521 141 559
rect 95 487 101 521
rect 135 487 141 521
rect 95 449 141 487
rect 95 415 101 449
rect 135 415 141 449
rect 95 377 141 415
rect 95 343 101 377
rect 135 343 141 377
rect 95 305 141 343
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -343 141 -305
rect 95 -377 101 -343
rect 135 -377 141 -343
rect 95 -415 141 -377
rect 95 -449 101 -415
rect 135 -449 141 -415
rect 95 -487 141 -449
rect 95 -521 101 -487
rect 135 -521 141 -487
rect 95 -559 141 -521
rect 95 -593 101 -559
rect 135 -593 141 -559
rect 95 -631 141 -593
rect 95 -665 101 -631
rect 135 -665 141 -631
rect 95 -703 141 -665
rect 95 -737 101 -703
rect 135 -737 141 -703
rect 95 -775 141 -737
rect 95 -809 101 -775
rect 135 -809 141 -775
rect 95 -847 141 -809
rect 95 -881 101 -847
rect 135 -881 141 -847
rect 95 -919 141 -881
rect 95 -953 101 -919
rect 135 -953 141 -919
rect 95 -991 141 -953
rect 95 -1025 101 -991
rect 135 -1025 141 -991
rect 95 -1063 141 -1025
rect 95 -1097 101 -1063
rect 135 -1097 141 -1063
rect 95 -1135 141 -1097
rect 95 -1169 101 -1135
rect 135 -1169 141 -1135
rect 95 -1207 141 -1169
rect 95 -1241 101 -1207
rect 135 -1241 141 -1207
rect 95 -1279 141 -1241
rect 95 -1313 101 -1279
rect 135 -1313 141 -1279
rect 95 -1351 141 -1313
rect 95 -1385 101 -1351
rect 135 -1385 141 -1351
rect 95 -1423 141 -1385
rect 95 -1457 101 -1423
rect 135 -1457 141 -1423
rect 95 -1500 141 -1457
rect -88 -1538 -30 -1532
rect -88 -1572 -76 -1538
rect -42 -1572 -30 -1538
rect -88 -1578 -30 -1572
rect 30 -1538 88 -1532
rect 30 -1572 42 -1538
rect 76 -1572 88 -1538
rect 30 -1578 88 -1572
<< properties >>
string FIXED_BBOX -232 -1657 232 1657
<< end >>
