magic
tech sky130A
magscale 1 1
timestamp 1737500400
<< checkpaint >>
rect 0 0 495 160
<< ndiff >>
rect 315 20 405 60
rect 315 60 405 100
rect 315 100 405 140
<< ptap >>
rect -45 -20 45 20
rect -45 20 45 60
rect -45 60 45 100
rect -45 100 45 140
rect -45 140 45 180
<< poly >>
rect 135 -8 435 8
rect 135 72 435 88
rect 135 152 435 168
rect 135 60 225 100
<< locali >>
rect 135 65 225 95
rect -45 -20 45 20
rect -45 20 45 60
rect 315 25 405 55
rect 315 25 405 55
rect -45 60 45 100
rect -45 60 45 100
rect 135 65 225 95
rect -45 100 45 140
rect 315 105 405 135
rect 315 105 405 135
rect -45 140 45 180
<< pcontact >>
rect 150 70 165 80
rect 150 80 165 90
rect 165 70 195 80
rect 165 80 195 90
rect 195 70 210 80
rect 195 80 210 90
<< ptapc >>
rect -15 20 15 60
rect -15 100 15 140
<< ndcontact >>
rect 330 30 345 40
rect 330 40 345 50
rect 345 30 375 40
rect 345 40 375 50
rect 375 30 390 40
rect 375 40 390 50
rect 330 110 345 120
rect 330 120 345 130
rect 345 110 375 120
rect 345 120 375 130
rect 375 110 390 120
rect 375 120 390 130
<< pwell >>
rect -75 -60 495 220
<< labels >>
flabel locali s 135 65 225 95 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 315 25 405 55 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -45 60 45 100 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 315 105 405 135 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 495 160
<< end >>
