magic
tech sky130A
magscale 1 1
timestamp 1737500400
<< checkpaint >>
rect 0 0 724 1720
<< locali >>
rect 8 8 716 64
rect 64 8 660 64
rect 8 8 716 64
rect 64 1656 660 1712
rect 8 1656 716 1712
rect 8 64 64 1656
rect 8 8 64 1712
rect 660 64 716 1656
rect 660 8 716 1712
rect 8 8 716 64
rect 398 1460 542 1580
rect 182 1460 326 1580
<< ptapc >>
rect 82 16 122 56
rect 122 16 162 56
rect 162 16 202 56
rect 202 16 242 56
rect 242 16 282 56
rect 282 16 322 56
rect 322 16 362 56
rect 362 16 402 56
rect 402 16 442 56
rect 442 16 482 56
rect 482 16 522 56
rect 522 16 562 56
rect 562 16 602 56
rect 602 16 642 56
rect 82 1664 122 1704
rect 122 1664 162 1704
rect 162 1664 202 1704
rect 202 1664 242 1704
rect 242 1664 282 1704
rect 282 1664 322 1704
rect 322 1664 362 1704
rect 362 1664 402 1704
rect 402 1664 442 1704
rect 442 1664 482 1704
rect 482 1664 522 1704
rect 522 1664 562 1704
rect 562 1664 602 1704
rect 602 1664 642 1704
rect 16 80 56 120
rect 16 120 56 160
rect 16 160 56 200
rect 16 200 56 240
rect 16 240 56 280
rect 16 280 56 320
rect 16 320 56 360
rect 16 360 56 400
rect 16 400 56 440
rect 16 440 56 480
rect 16 480 56 520
rect 16 520 56 560
rect 16 560 56 600
rect 16 600 56 640
rect 16 640 56 680
rect 16 680 56 720
rect 16 720 56 760
rect 16 760 56 800
rect 16 800 56 840
rect 16 840 56 880
rect 16 880 56 920
rect 16 920 56 960
rect 16 960 56 1000
rect 16 1000 56 1040
rect 16 1040 56 1080
rect 16 1080 56 1120
rect 16 1120 56 1160
rect 16 1160 56 1200
rect 16 1200 56 1240
rect 16 1240 56 1280
rect 16 1280 56 1320
rect 16 1320 56 1360
rect 16 1360 56 1400
rect 16 1400 56 1440
rect 16 1440 56 1480
rect 16 1480 56 1520
rect 16 1520 56 1560
rect 16 1560 56 1600
rect 16 1600 56 1640
rect 668 80 708 120
rect 668 120 708 160
rect 668 160 708 200
rect 668 200 708 240
rect 668 240 708 280
rect 668 280 708 320
rect 668 320 708 360
rect 668 360 708 400
rect 668 400 708 440
rect 668 440 708 480
rect 668 480 708 520
rect 668 520 708 560
rect 668 560 708 600
rect 668 600 708 640
rect 668 640 708 680
rect 668 680 708 720
rect 668 720 708 760
rect 668 760 708 800
rect 668 800 708 840
rect 668 840 708 880
rect 668 880 708 920
rect 668 920 708 960
rect 668 960 708 1000
rect 668 1000 708 1040
rect 668 1040 708 1080
rect 668 1080 708 1120
rect 668 1120 708 1160
rect 668 1160 708 1200
rect 668 1200 708 1240
rect 668 1240 708 1280
rect 668 1280 708 1320
rect 668 1320 708 1360
rect 668 1360 708 1400
rect 668 1400 708 1440
rect 668 1440 708 1480
rect 668 1480 708 1520
rect 668 1520 708 1560
rect 668 1560 708 1600
rect 668 1600 708 1640
<< ptap >>
rect 0 0 724 72
rect 0 1648 724 1720
rect 0 0 72 1720
rect 652 0 724 1720
use JNWTR_RES2 XA1 
transform 1 0 200 0 1 200
box 200 200 524 1520
<< labels >>
flabel locali s 8 8 716 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 398 1460 542 1580 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 182 1460 326 1580 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 724 1720
<< end >>
