
*.subckt CAPX1 A B
*C1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
*.ends


.subckt CAPX4 A B
XA1 A B CAPX1 xoffset=8 yoffset=0
XA2 A B CAPX1 yoffset=6
XB1 A B CAPX1 xoffset=8
XB2 A B CAPX1 yoffset=6
.ends
