magic
tech sky130A
magscale 1 1
timestamp 1737500400
<< checkpaint >>
rect 0 0 495 160
<< pdiff >>
rect 90 20 180 60
rect 90 60 180 100
rect 90 100 180 140
<< ntap >>
rect 450 -20 540 20
rect 450 20 540 60
rect 450 60 540 100
rect 450 100 540 140
rect 450 140 540 180
<< poly >>
rect 60 -8 360 8
rect 60 72 360 88
rect 60 152 360 168
rect 270 60 360 100
<< locali >>
rect 270 65 360 95
rect 450 -20 540 20
rect 90 25 180 55
rect 90 25 180 55
rect 450 20 540 60
rect 270 65 360 95
rect 450 60 540 100
rect 450 60 540 100
rect 90 105 180 135
rect 90 105 180 135
rect 450 100 540 140
rect 450 140 540 180
<< pcontact >>
rect 285 70 300 80
rect 285 80 300 90
rect 300 70 330 80
rect 300 80 330 90
rect 330 70 345 80
rect 330 80 345 90
<< ntapc >>
rect 480 20 510 60
rect 480 100 510 140
<< pdcontact >>
rect 105 30 120 40
rect 105 40 120 50
rect 120 30 150 40
rect 120 40 150 50
rect 150 30 165 40
rect 150 40 165 50
rect 105 110 120 120
rect 105 120 120 130
rect 120 110 150 120
rect 120 120 150 130
rect 150 110 165 120
rect 150 120 165 130
<< nwell >>
rect 0 -60 570 220
<< labels >>
flabel locali s 270 65 360 95 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 90 25 180 55 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 450 60 540 100 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 90 105 180 135 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 495 160
<< end >>
