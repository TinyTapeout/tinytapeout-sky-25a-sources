* NGSPICE file created from tt_um_13hihi31_tdc_parax.ext - technology: sky130A

.subckt tt_um_13hihi31_tdc_parax clk ena rst_n ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[1] ui_in[5]
+ uo_out[7] ui_in[7] uio_in[0] uo_out[6] ui_in[4] uo_out[5] ua[0] uo_out[4] uo_out[0]
+ ui_in[3] uo_out[3] ui_in[6] ui_in[2] ui_in[1] uio_in[6] VGND VDPWR ui_in[0] uo_out[2]
X0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 VDPWR.t294 VDPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1 tdc_0.start_buffer_0.start_delay.t7 tdc_0.start_buffer_0.start_buff.t10 VDPWR.t326 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X2 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VDPWR.t427 VDPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X3 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X4 tdc_0.vernier_delay_line_0.stop_strong.t15 a_9330_16954.t8 VGND.t561 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5 a_10958_39338.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 a_10108_39954.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X6 a_10108_28544.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X7 VDPWR.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30598# VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X8 VGND.t1 input_stage_andpwr_0.fine_delay_unit_0.in a_24790_6936# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X9 a_10958_23364.t7 tdc_0.vernier_delay_line_0.stop_strong.t32 VGND.t453 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X10 a_24240_11366# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VDPWR.t560 VDPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 a_13254_26412# VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X12 tdc_0.vernier_delay_line_0.stop_strong.t31 a_9330_16954.t9 VDPWR.t607 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X13 a_10108_35390.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 a_13254_35540# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X15 VDPWR.t360 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X16 VGND.t290 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 a_25060_21092# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X17 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 a_10958_39338.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X18 VDPWR.t149 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 a_24240_26106# VDPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X19 a_10958_37056.t8 tdc_0.vernier_delay_line_0.stop_strong.t33 VGND.t161 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X20 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 a_10108_26262.t2 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X21 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 VDPWR.t465 VDPWR.t467 VDPWR.t466 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X22 VGND.t162 tdc_0.vernier_delay_line_0.stop_strong.t34 a_10958_23364.t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X23 a_9330_14344# a_9330_14054# VGND.t554 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X24 uo_out[6].t0 a_12310_37398# VGND.t226 VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X25 VGND.t93 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 VGND.t203 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X27 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 a_10108_35390.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X28 a_9330_16954.t3 a_9330_15794# VGND.t528 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X29 VDPWR.t221 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 a_24240_23158# VDPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X30 a_7140_10670# variable_delay_dummy_0.out VDPWR.t469 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X31 variable_delay_short_0.in a_23820_8460# VGND.t207 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X32 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 VGND.t291 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X33 VGND.t289 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X34 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 VDPWR.t413 VDPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X35 VDPWR.t540 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 VDPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X36 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 a_10958_39338.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X37 a_10958_37056.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 a_10108_37144# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X38 VGND.t227 tdc_0.vernier_delay_line_0.stop_strong.t35 a_10958_34774.t8 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X39 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 VDPWR.t542 VDPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X40 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12308_33296# a_12420_33258# VDPWR.t264 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X41 VGND.t269 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X42 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VGND.t303 VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X43 a_13254_35162# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 uo_out[5].t1 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X44 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 VDPWR.t296 VDPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X45 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 VGND.t143 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X46 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 ui_in[5].t0 VDPWR.t553 VDPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X47 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 VDPWR.t306 VDPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X48 VGND.t559 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 a_12310_25988# VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X49 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12308_40142# a_12420_40104# VDPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X50 a_10108_28544.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 a_10958_27928.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X51 tdc_0.start_buffer_0.start_buff.t3 a_7140_10670# VGND.t150 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X52 VDPWR.t242 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 a_24240_17262# VDPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X53 VGND.t250 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 VGND.t249 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X54 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND.t359 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X55 VGND.t115 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 a_12310_32834# VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X56 a_16292_6966# input_stage_0.fine_delay_unit_0.in a_16292_6702# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X57 VDPWR.t502 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 a_15680_14582# VDPWR.t501 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X58 a_10108_35390.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 a_10958_34774.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X59 a_10108_30826.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X60 a_9330_15794# a_9330_15504# VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X61 VDPWR.t362 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X62 VDPWR.t411 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 VDPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X63 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 VGND.t307 VGND.t306 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X64 VGND.t224 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 a_25060_18144# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X65 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 VGND.t501 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 VDPWR.t308 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 VDPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X67 a_10108_28544.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 a_10958_27928.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X68 a_24790_8050# input_stage_andpwr_0.fine_delay_unit_1.in a_23820_8460# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X69 tdc_0.vernier_delay_line_0.stop_strong.t30 a_9330_16954.t10 VDPWR.t608 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X70 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 VDPWR.t615 VGND.t410 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X71 uo_out[0].t0 a_12310_23706# VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X72 a_10958_25646.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 a_10108_26262.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X73 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 VDPWR.t244 VDPWR.t243 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X74 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VDPWR.t383 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X75 a_25060_26988# VGND.t17 variable_delay_short_0.variable_delay_unit_5.out VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X76 VDPWR.t423 tdc_0.start_buffer_0.start_buff.t11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 VDPWR.t422 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X77 tdc_0.vernier_delay_line_0.stop_strong.t29 a_9330_16954.t11 VDPWR.t609 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X78 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VDPWR.t504 VDPWR.t503 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X79 a_10958_34774.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 a_10108_35390.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X80 uo_out[3].t2 a_12310_30552# VGND.t553 VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X81 VGND.t100 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 a_16500_12516# VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X82 VGND.t480 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 VGND.t479 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X83 VGND.t228 tdc_0.vernier_delay_line_0.stop_strong.t36 a_10958_32492.t9 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X84 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VDPWR.t407 VDPWR.t406 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X85 VGND.t475 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 a_25060_26988# VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X86 VDPWR.t531 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 VDPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X87 VGND.t109 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X88 a_10958_23364.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 a_10108_23452# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X89 VGND.t537 input_stage_0.fine_delay_unit_1.in a_16292_8344# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X90 VGND.t159 tdc_0.vernier_delay_line_0.stop_strong.t37 a_10958_39338.t7 VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X91 a_23820_7082# input_stage_andpwr_0.fine_delay_unit_0.in a_24790_6672# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X92 VDPWR.t127 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 VDPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X93 VDPWR.t278 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 VDPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X94 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X95 VGND.t160 tdc_0.vernier_delay_line_0.stop_strong.t38 a_10958_25646.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X96 VGND.t507 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 VGND.t506 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X97 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 ui_in[5].t1 VGND.t524 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X98 VDPWR.t353 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 VDPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X99 tdc_0.vernier_delay_line_0.stop_strong.t14 a_9330_16954.t12 VGND.t131 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X100 VDPWR.t532 tdc_0.vernier_delay_line_0.stop_strong.t39 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X101 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 VDPWR.t88 VDPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X102 a_10958_34774.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 a_10108_35390.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X103 a_13254_30598# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 uo_out[3].t0 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X104 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 VDPWR.t314 VDPWR.t313 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X105 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 VGND.t279 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X106 VGND.t490 tdc_0.vernier_delay_line_0.stop_strong.t40 a_10958_32492.t8 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X107 variable_delay_short_0.variable_delay_unit_5.forward.t1 variable_delay_short_0.variable_delay_unit_5.in.t2 VDPWR.t579 VDPWR.t466 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X108 a_9330_14344# a_9330_14054# VDPWR.t597 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X109 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 VGND.t434 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X110 a_16292_8080# input_stage_0.fine_delay_unit_1.in a_15322_8490# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X111 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 tdc_0.start_buffer_0.start_buff.t12 VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X112 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 a_10958_25646.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X113 a_24790_6672# input_stage_andpwr_0.fine_delay_unit_0.in a_23820_7082# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X114 a_9330_16954.t7 a_9330_15794# VDPWR.t557 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X115 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 VDPWR.t344 VDPWR.t343 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X116 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VDPWR.t550 VDPWR.t549 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X117 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VDPWR.t616 VGND.t409 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X118 a_10958_23364.t5 tdc_0.vernier_delay_line_0.stop_strong.t41 VGND.t325 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X119 a_10108_30826.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 a_10958_30210.t8 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X120 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 VGND.t179 VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X121 a_25060_20210# ui_in[5].t2 VGND.t261 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X122 a_10958_30210.t4 tdc_0.vernier_delay_line_0.stop_strong.t42 VGND.t326 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X123 a_10108_23980.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 a_10958_23364.t9 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X124 variable_delay_short_0.variable_delay_unit_4.in.t1 variable_delay_short_0.variable_delay_unit_3.in.t2 VDPWR.t251 VDPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X125 VDPWR.t415 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 VDPWR.t414 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X126 a_15322_8490# input_stage_0.fine_delay_unit_1.in a_16292_8080# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X127 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 VGND.t305 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X128 a_10958_39338.t6 tdc_0.vernier_delay_line_0.stop_strong.t43 VGND.t512 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X129 VDPWR.t517 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 VDPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X130 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 tdc_0.start_buffer_0.start_delay.t8 VDPWR.t506 VDPWR.t505 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X131 VDPWR.t286 ui_in[5].t3 a_24240_21092# VDPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X132 a_13254_24130# uo_out[0].t4 VGND.t342 VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X133 VGND.t360 ui_in[5].t4 a_25060_20210# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X134 VGND.t301 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X135 a_13254_33258# uo_out[4].t4 VGND.t484 VGND.t483 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X136 VGND.t513 tdc_0.vernier_delay_line_0.stop_strong.t44 a_10958_30210.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X137 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND.t503 VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X138 a_24240_24040# ui_in[4].t0 VDPWR.t98 VDPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X139 VGND.t523 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X140 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 a_10958_34774.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X141 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 VDPWR.t527 VDPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X142 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 VDPWR.t524 VDPWR.t523 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X143 a_13254_40104# uo_out[7].t4 VGND.t202 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X144 variable_delay_short_0.variable_delay_unit_5.forward.t0 variable_delay_short_0.variable_delay_unit_5.in.t3 VGND.t192 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X145 a_9330_15214# a_9330_14924# VGND.t94 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X146 a_24240_21092# ui_in[5].t5 VDPWR.t417 VDPWR.t416 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X147 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VDPWR.t62 VDPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X148 VDPWR.t143 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28316# VDPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X149 VGND.t102 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X150 a_25060_18144# variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X151 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 VGND.t275 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X152 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 VDPWR.t429 VDPWR.t428 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X153 tdc_0.vernier_delay_line_0.stop_strong.t13 a_9330_16954.t13 VGND.t132 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X154 tdc_0.vernier_delay_line_0.start_pos.t5 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 VDPWR.t575 VDPWR.t574 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X155 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12308_37860# a_12420_37822# VDPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X156 VGND.t152 ui_in[7].t0 a_25060_14314# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X157 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 a_13254_30976# VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X158 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 VGND.t182 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X159 tdc_0.vernier_delay_line_0.stop_strong.t12 a_9330_16954.t14 VGND.t133 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X160 VDPWR.t321 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X161 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X162 a_24240_18144# ui_in[6].t0 VDPWR.t591 VDPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X163 tdc_0.vernier_delay_line_0.stop_strong.t11 a_9330_16954.t15 VGND.t106 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X164 a_25284_5108# uio_in[6].t0 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X165 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t219 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X166 VDPWR.t323 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VDPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X167 VGND.t308 uio_in[0].t0 a_25060_11366# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X168 variable_delay_short_0.variable_delay_unit_4.in.t0 variable_delay_short_0.variable_delay_unit_3.in.t3 VGND.t481 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X169 VDPWR.t409 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VDPWR.t408 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X170 VGND.t469 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X171 tdc_0.vernier_delay_line_0.stop_strong.t28 a_9330_16954.t16 VDPWR.t110 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X172 tdc_0.vernier_delay_line_0.start_neg.t7 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X173 a_24240_15196# ui_in[7].t1 VDPWR.t166 VDPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X174 VGND.t277 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X175 VDPWR.t370 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VDPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X176 VDPWR.t564 tdc_0.vernier_delay_line_0.start_pos.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 VDPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X177 VGND.t36 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_13254_39726# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X178 a_15680_12516# VDPWR.t462 VDPWR.t464 VDPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X179 VGND.t373 tdc_0.start_buffer_0.start_delay.t9 tdc_0.start_buffer_0.start_buff.t9 VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X180 VDPWR.t68 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VDPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X181 a_10108_33108.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 a_10958_32492.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X182 VDPWR.t593 ui_in[6].t1 a_24240_18144# VDPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X183 a_25060_26106# VDPWR.t617 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X184 VDPWR.t300 tdc_0.start_buffer_0.start_buff.t13 tdc_0.start_buffer_0.start_delay.t6 VDPWR.t299 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X185 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 variable_delay_dummy_0.variable_delay_unit_1.in.t2 VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X186 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X187 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t320 VDPWR.t319 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X188 a_9330_13764# variable_delay_short_0.out VGND.t127 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X189 VDPWR.t461 VDPWR.t459 a_15680_15464# VDPWR.t460 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X190 VGND.t234 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X191 VGND.t78 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X192 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 VDPWR.t614 VDPWR.t613 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X193 a_24240_26988# VGND.t562 variable_delay_short_0.variable_delay_unit_5.out VDPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X194 VDPWR.t124 tdc_0.vernier_delay_line_0.stop_strong.t45 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VDPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X195 a_25060_23158# ui_in[4].t1 VGND.t91 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X196 VDPWR.t270 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 VDPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X197 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t398 VDPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X198 VGND.t184 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X199 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VDPWR.t80 VDPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X200 VDPWR.t458 VDPWR.t456 a_24240_26988# VDPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X201 VDPWR.t181 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 VDPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X202 a_10958_30210.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 a_10108_30826.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X203 tdc_0.start_buffer_0.start_buff.t7 a_7140_10670# VDPWR.t162 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X204 a_23820_7082# input_stage_andpwr_0.fine_delay_unit_0.in VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X205 a_16786_5138# uio_in[6].t1 VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X206 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 VDPWR.t349 VDPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X207 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.start_pos.t9 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X208 VDPWR.t500 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37444# VDPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X209 a_24790_8314# ui_in[2].t0 a_24790_8050# VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X210 VDPWR.t17 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X211 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X212 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 VGND.t51 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X213 tdc_0.start_buffer_0.start_buff.t2 a_7140_10670# VGND.t149 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X214 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VGND.t73 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X215 VDPWR.t475 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 VDPWR.t474 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X216 VDPWR.t371 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X217 tdc_0.start_buffer_0.start_delay.t1 tdc_0.start_buffer_0.start_buff.t14 VGND.t382 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X218 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VDPWR.t133 VDPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X219 a_12420_26412# uo_out[1].t4 VDPWR.t263 VDPWR.t262 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X220 a_9330_15214# a_9330_14924# VDPWR.t103 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X221 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 VGND.t248 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X222 VGND.t85 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X223 tdc_0.vernier_delay_line_0.start_pos.t2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X224 VGND.t49 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X225 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 tdc_0.vernier_delay_line_0.start_neg.t8 VDPWR.t342 VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X226 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 VDPWR.t334 VDPWR.t333 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X227 tdc_0.vernier_delay_line_0.stop_strong.t27 a_9330_16954.t17 VDPWR.t111 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X228 VDPWR.t42 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 VDPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X229 a_15322_8490# input_stage_0.fine_delay_unit_1.in VDPWR.t573 VDPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X230 VGND.t45 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X231 VGND.t116 tdc_0.vernier_delay_line_0.stop_strong.t46 a_10958_37056.t7 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X232 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 a_10958_30210.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X233 tdc_0.vernier_delay_line_0.stop_strong.t26 a_9330_16954.t18 VDPWR.t172 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X234 tdc_0.vernier_delay_line_0.start_neg.t4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X235 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 VDPWR.t604 VDPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X236 VDPWR.t325 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 a_12310_28270# VDPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X237 variable_delay_dummy_0.in a_15322_8490# VDPWR.t78 VDPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X238 VGND.t406 VDPWR.t618 a_16500_14582# VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X239 tdc_0.vernier_delay_line_0.stop_strong.t25 a_9330_16954.t19 VDPWR.t173 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X240 a_12420_32880# a_12310_32834# uo_out[4].t1 VDPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X241 VGND.t198 tdc_0.vernier_delay_line_0.stop_strong.t47 a_10958_27928.t8 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X242 VGND.t12 tdc_0.vernier_delay_line_0.start_pos.t10 tdc_0.vernier_delay_line_0.start_neg.t0 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X243 VDPWR.t168 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 a_12310_37398# VDPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X244 a_13254_28316# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 uo_out[2].t0 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X245 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t48 VDPWR.t215 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X246 a_16292_8344# uio_in[3].t0 a_16292_8080# VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X247 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X248 a_24790_6936# ui_in[0].t0 a_24790_6672# VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X249 VDPWR.t336 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 a_24240_20210# VDPWR.t335 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X250 a_13254_37822# uo_out[6].t4 VGND.t460 VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X251 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out VDPWR.t332 VDPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X252 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t49 VDPWR.t216 VDPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X253 VDPWR.t392 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_23752# VDPWR.t391 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X254 a_16500_14582# VDPWR.t619 VGND.t404 VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X255 VDPWR.t566 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_32880# VDPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X256 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 a_13254_28694# VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X257 a_10958_25646.t10 tdc_0.vernier_delay_line_0.stop_strong.t50 VGND.t199 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X258 VGND.t452 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 a_12310_39680# VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X259 VDPWR.t70 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VDPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X260 a_9330_13764# variable_delay_short_0.out VDPWR.t141 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X261 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 a_10108_39426# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X262 uo_out[5].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t400 VDPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X263 VGND.t195 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26034# VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X264 VDPWR.t72 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X265 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 ui_in[6].t2 VDPWR.t567 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X266 a_10108_37672.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X267 a_24240_18144# variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out VDPWR.t558 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X268 VDPWR.t123 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X269 VDPWR.t131 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 a_24240_14314# VDPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X270 a_15680_15464# VGND.t563 variable_delay_dummy_0.variable_delay_unit_1.out VDPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X271 a_25060_12248# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND.t529 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X272 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 ui_in[7].t2 VDPWR.t137 VDPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X273 a_12420_26034# a_12310_25988# uo_out[1].t1 VDPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X274 VGND.t189 tdc_0.vernier_delay_line_0.start_neg.t9 tdc_0.vernier_delay_line_0.start_pos.t6 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X275 VDPWR.t23 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 a_15680_11634# VDPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X276 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 a_10108_28544.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X277 uo_out[7].t2 a_12310_39680# VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X278 a_12420_35540# uo_out[5].t4 VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X279 VDPWR.t562 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 a_24240_11366# VDPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X280 VDPWR.t536 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VDPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X281 VGND.t390 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X282 VGND.t246 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X283 VDPWR.t292 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VDPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X284 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X285 VGND.t464 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 tdc_0.vernier_delay_line_0.start_pos.t1 VGND.t463 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X286 VDPWR.t600 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 a_12310_23706# VDPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X287 a_10958_39338.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 a_10108_39426# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X288 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.start_neg.t10 VGND.t364 VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X289 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 VDPWR.t513 VDPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X290 VGND.t259 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X291 VDPWR.t156 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 a_12310_30552# VDPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X292 tdc_0.vernier_delay_line_0.stop_strong.t10 a_9330_16954.t20 VGND.t163 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X293 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VGND.t466 VGND.t465 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X294 VDPWR.t544 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 VDPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X295 VGND.t204 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 a_25060_24040# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X296 a_13254_37444# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 uo_out[6].t3 VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X297 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 VDPWR.t207 VDPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X298 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VGND.t191 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X299 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 VDPWR.t351 VDPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X300 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 a_10108_25734# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X301 VGND.t478 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 a_25060_21092# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X302 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 VGND.t344 VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X303 a_10108_23980.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X304 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 ui_in[6].t3 VGND.t534 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X305 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 VDPWR.t117 VDPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X306 a_10958_39338.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 a_10108_39426# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X307 a_10108_37672.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 a_10958_37056.t9 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X308 VGND.t171 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 a_12310_35116# VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X309 variable_delay_short_0.variable_delay_unit_5.in.t1 variable_delay_short_0.variable_delay_unit_4.in.t2 VDPWR.t368 VDPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X310 a_10958_34774.t7 tdc_0.vernier_delay_line_0.stop_strong.t51 VGND.t337 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X311 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 VGND.t267 VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X312 VDPWR.t236 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VDPWR.t235 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X313 input_stage_0.fine_delay_unit_1.in a_15322_7112# VDPWR.t473 VDPWR.t472 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X314 VGND.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35162# VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X315 input_stage_andpwr_0.fine_delay_unit_1.in a_23820_7082# VGND.t166 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X316 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 ui_in[7].t3 VGND.t125 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X317 tdc_0.vernier_delay_line_0.stop_strong.t9 a_9330_16954.t21 VGND.t355 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X318 VDPWR.t96 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 VDPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X319 a_10958_27928.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 a_10108_28544.t5 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X320 uo_out[1].t0 a_12310_25988# VGND.t43 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X321 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VDPWR.t620 VGND.t402 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X322 VDPWR.t170 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X323 tdc_0.vernier_delay_line_0.stop_strong.t8 a_9330_16954.t22 VGND.t356 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X324 VDPWR.t56 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 VDPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X325 a_10108_37672.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 a_10958_37056.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X326 a_12420_30976# uo_out[3].t4 VDPWR.t382 VDPWR.t381 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X327 input_stage_andpwr_0.nand_gate_0.out uio_in[6].t2 ua[0].t1 ua[0].t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X328 VGND.t358 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 a_25060_15196# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X329 uo_out[4].t0 a_12310_32834# VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X330 VGND.t265 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X331 VDPWR.t121 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 VDPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X332 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 a_10108_30826.t4 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X333 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 a_10958_27928.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X334 variable_delay_short_0.variable_delay_unit_3.in.t1 variable_delay_short_0.variable_delay_unit_2.in.t2 VDPWR.t387 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X335 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t185 VDPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X336 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 VDPWR.t304 VDPWR.t303 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X337 a_10958_27928.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 a_10108_28544.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X338 a_24790_8314# input_stage_andpwr_0.fine_delay_unit_1.in a_24790_8050# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X339 a_13254_23752# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 uo_out[0].t2 VGND.t253 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X340 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t385 VDPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X341 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VDPWR.t255 VDPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X342 VGND.t333 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X343 a_10958_32492.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 a_10108_32580# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X344 variable_delay_short_0.variable_delay_unit_2.in.t0 variable_delay_short_0.variable_delay_unit_1.in.t2 VDPWR.t605 VDPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X345 a_10958_37056.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 a_10108_37672.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X346 a_16292_6702# input_stage_0.fine_delay_unit_0.in a_15322_7112# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X347 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 tdc_0.start_buffer_0.start_buff.t15 VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X348 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward.t2 a_15680_14582# VDPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X349 a_9330_14634# a_9330_14344# VGND.t244 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X350 VGND.t338 tdc_0.vernier_delay_line_0.stop_strong.t52 a_10958_34774.t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X351 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VDPWR.t453 VDPWR.t455 VDPWR.t454 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X352 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X353 a_16500_12516# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X354 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 a_13254_24130# VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X355 a_10958_25646.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 a_10108_25734# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X356 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 VDPWR.t375 VDPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X357 a_10108_23980.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 a_10958_23364.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X358 a_9330_16954.t2 a_9330_15794# VGND.t527 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X359 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X360 a_10108_33108.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X361 tdc_0.start_buffer_0.start_buff.t6 a_7140_10670# VDPWR.t161 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X362 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 a_10958_27928.t2 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X363 VGND.t505 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 a_16500_15464# VGND.t504 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X364 variable_delay_short_0.variable_delay_unit_5.in.t0 variable_delay_short_0.variable_delay_unit_4.in.t3 VGND.t241 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X365 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 a_10108_34862# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X366 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 VGND.t113 VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X367 tdc_0.start_buffer_0.start_delay.t5 tdc_0.start_buffer_0.start_buff.t16 VDPWR.t198 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X368 a_25060_15196# variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_1.out VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X369 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 VDPWR.t481 VDPWR.t480 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X370 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 a_10958_34774.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X371 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 a_10108_23980.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X372 input_stage_0.nand_gate_0.out uio_in[6].t3 VDPWR.t140 VDPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X373 a_10958_32492.t7 tdc_0.vernier_delay_line_0.stop_strong.t53 VGND.t229 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X374 VGND.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30598# VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X375 tdc_0.vernier_delay_line_0.stop_strong.t24 a_9330_16954.t23 VDPWR.t405 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X376 VGND.t31 input_stage_0.fine_delay_unit_0.in a_16292_6966# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X377 a_25060_12248# variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X378 tdc_0.start_buffer_0.start_buff.t1 a_7140_10670# VGND.t148 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X379 VGND.t539 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X380 VDPWR.t272 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 VDPWR.t271 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X381 a_10958_25646.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 a_10108_25734# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X382 a_24790_6936# input_stage_andpwr_0.fine_delay_unit_0.in a_24790_6672# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X383 VGND.t139 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X384 VDPWR.t552 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 VDPWR.t551 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X385 VGND.t230 tdc_0.vernier_delay_line_0.stop_strong.t54 a_10958_23364.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X386 variable_delay_short_0.variable_delay_unit_3.in.t0 variable_delay_short_0.variable_delay_unit_2.in.t3 VGND.t130 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X387 a_25060_24040# variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.out VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X388 VGND.t509 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VGND.t508 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X389 a_10958_30210.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 a_10108_30826.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X390 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X391 a_24240_12248# uio_in[0].t1 VDPWR.t355 VDPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X392 a_12420_39726# a_12310_39680# uo_out[7].t3 VDPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X393 VGND.t477 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 a_25060_26988# VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X394 VDPWR.t519 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 VDPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X395 variable_delay_short_0.variable_delay_unit_2.in.t1 variable_delay_short_0.variable_delay_unit_1.in.t3 VGND.t560 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X396 a_10958_23364.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 a_10108_23980.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X397 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 VDPWR.t90 VDPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X398 tdc_0.vernier_delay_line_0.stop_strong.t23 a_9330_16954.t24 VDPWR.t192 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X399 a_16292_8080# input_stage_0.fine_delay_unit_1.in a_15322_8490# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X400 VGND.t547 tdc_0.vernier_delay_line_0.stop_strong.t55 a_10958_39338.t5 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X401 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 VGND.t541 VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X402 variable_delay_dummy_0.variable_delay_unit_1.in.t0 variable_delay_dummy_0.in VGND.t426 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X403 tdc_0.vernier_delay_line_0.stop_strong.t22 a_9330_16954.t25 VDPWR.t193 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X404 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.stop_strong.t56 VDPWR.t588 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X405 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 VDPWR.t195 VDPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X406 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X407 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 VDPWR.t74 VDPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X408 a_25060_20210# ui_in[5].t6 VGND.t361 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X409 a_10108_33108.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 a_10958_32492.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X410 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 a_13254_33258# VGND.t221 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X411 a_10958_30210.t2 tdc_0.vernier_delay_line_0.stop_strong.t57 VGND.t235 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X412 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 VGND.t252 VGND.t251 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X413 VDPWR.t611 ui_in[4].t2 a_24240_24040# VDPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X414 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 VGND.t521 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X415 a_10958_34774.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 a_10108_34862# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X416 VDPWR.t529 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 VDPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X417 VDPWR.t92 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 VDPWR.t91 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X418 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 tdc_0.start_buffer_0.start_buff.t17 VGND.t381 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X419 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t316 VDPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X420 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 a_13254_40104# VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X421 a_10958_23364.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 a_10108_23980.t2 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X422 VDPWR.t230 tdc_0.start_buffer_0.start_delay.t10 tdc_0.start_buffer_0.start_buff.t8 VDPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X423 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 VGND.t197 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X424 VDPWR.t302 ui_in[5].t7 a_24240_21092# VDPWR.t301 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X425 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t479 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X426 VGND.t260 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 a_25060_18144# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X427 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 variable_delay_dummy_0.variable_delay_unit_1.in.t3 VDPWR.t598 VDPWR.t454 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X428 a_9330_14634# a_9330_14344# VDPWR.t265 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X429 a_24790_8050# input_stage_andpwr_0.fine_delay_unit_1.in a_23820_8460# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X430 a_25060_14314# ui_in[7].t4 VGND.t151 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X431 VDPWR.t257 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 VDPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X432 VGND.t88 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X433 VDPWR.t58 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 VDPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X434 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X435 VGND.t319 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X436 a_9330_16954.t6 a_9330_15794# VDPWR.t556 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X437 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 a_10108_39954.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X438 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 a_10958_37056.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X439 input_stage_andpwr_0.nand_gate_0.out VDPWR.t621 a_25284_5108# VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X440 VDPWR.t258 tdc_0.vernier_delay_line_0.stop_strong.t58 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X441 VGND.t455 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 VGND.t454 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X442 a_25060_11366# uio_in[0].t2 VGND.t299 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X443 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_3.in.t4 a_25060_17262# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X444 VDPWR.t240 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 VDPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X445 VGND.t420 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X446 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VGND.t489 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X447 VDPWR.t525 tdc_0.vernier_delay_line_0.stop_strong.t59 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X448 VDPWR.t164 ui_in[7].t5 a_24240_15196# VDPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X449 a_23820_8460# input_stage_andpwr_0.fine_delay_unit_1.in a_24790_8050# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X450 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in.t4 a_25060_14314# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X451 a_16500_15464# VGND.t15 variable_delay_dummy_0.variable_delay_unit_1.out VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X452 VGND.t545 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X453 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.start_pos.t11 VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X454 VDPWR.t452 VDPWR.t450 a_15680_12516# VDPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X455 a_10958_32492.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 a_10108_33108.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X456 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 VDPWR.t60 VDPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X457 VGND.t401 VDPWR.t622 a_16500_11634# VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X458 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 tdc_0.start_buffer_0.start_delay.t11 VGND.t371 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X459 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 VDPWR.t282 VDPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X460 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward.t2 a_25060_26106# VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X461 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 VDPWR.t232 VDPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X462 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 a_10108_30298# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X463 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VGND.t448 VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X464 uo_out[2].t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X465 tdc_0.vernier_delay_line_0.stop_strong.t7 a_9330_16954.t26 VGND.t180 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X466 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 VDPWR.t546 VDPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X467 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 VGND.t53 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X468 VDPWR.t496 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VDPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X469 VGND.t369 tdc_0.start_buffer_0.start_delay.t12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 VGND.t368 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X470 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 a_10958_30210.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X471 VDPWR.t38 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 VDPWR.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X472 tdc_0.vernier_delay_line_0.start_pos.t4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 VDPWR.t359 VDPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X473 a_10108_35390.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 a_10958_34774.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X474 VDPWR.t36 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 VDPWR.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X475 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t187 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X476 a_12420_28694# uo_out[2].t4 VDPWR.t105 VDPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X477 VGND.t450 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X478 VGND.t494 ui_in[3].t0 a_24790_8314# VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X479 tdc_0.vernier_delay_line_0.start_neg.t6 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X480 VGND.t111 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X481 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 a_10958_23364.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X482 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_1.out VDPWR.t509 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X483 VGND.t310 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X484 a_10958_39338.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 a_10108_39954.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X485 VDPWR.t5 tdc_0.vernier_delay_line_0.start_pos.t12 tdc_0.vernier_delay_line_0.start_neg.t1 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X486 a_15680_12516# variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out VDPWR.t511 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X487 a_16292_6966# uio_in[1].t0 a_16292_6702# VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X488 VGND.t315 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 VGND.t314 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X489 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 VDPWR.t477 VDPWR.t476 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X490 a_10958_30210.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 a_10108_30298# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X491 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 uio_in[0].t3 VDPWR.t340 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X492 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t64 VDPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X493 a_25060_26106# VDPWR.t623 VGND.t400 VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X494 a_24240_12248# variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out VDPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X495 VGND.t218 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X496 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12308_26450# a_12420_26412# VDPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X497 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 ui_in[4].t3 VDPWR.t612 VDPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X498 a_24240_24040# variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.out VDPWR.t3 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X499 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 VGND.t462 VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X500 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 VGND.t214 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X501 a_25060_23158# ui_in[4].t4 VGND.t222 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X502 VGND.t485 tdc_0.vernier_delay_line_0.stop_strong.t60 a_10958_37056.t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X503 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t61 VDPWR.t492 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X504 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12308_35578# a_12420_35540# VDPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X505 VDPWR.t449 VDPWR.t447 a_24240_26988# VDPWR.t448 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X506 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 VGND.t531 VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X507 a_10958_30210.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 a_10108_30298# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X508 VGND.t24 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 tdc_0.vernier_delay_line_0.start_neg.t3 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X509 a_9330_14054# a_9330_13764# VGND.t86 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X510 a_10958_27928.t7 tdc_0.vernier_delay_line_0.stop_strong.t62 VGND.t456 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X511 VDPWR.t425 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VDPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X512 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.start_pos.t13 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X513 uo_out[6].t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t581 VDPWR.t580 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X514 VGND.t129 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28316# VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X515 input_stage_andpwr_0.fine_delay_unit_0.in input_stage_andpwr_0.nand_gate_0.out VGND.t297 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X516 a_9330_15504# a_9330_15214# VGND.t425 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X517 a_10108_39954.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X518 VGND.t493 uio_in[4].t0 a_16292_8344# VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X519 VDPWR.t225 tdc_0.vernier_delay_line_0.start_neg.t11 tdc_0.vernier_delay_line_0.start_pos.t7 VDPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X520 a_9330_16954.t1 a_9330_15794# VGND.t526 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X521 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 VDPWR.t515 VDPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X522 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 a_13254_37822# VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X523 a_25060_17262# ui_in[6].t4 VGND.t298 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X524 tdc_0.vernier_delay_line_0.stop_strong.t6 a_9330_16954.t27 VGND.t136 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X525 VDPWR.t484 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 VDPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X526 tdc_0.start_buffer_0.start_buff.t5 a_7140_10670# VDPWR.t160 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X527 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward.t3 a_16500_14582# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X528 VGND.t59 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X529 tdc_0.vernier_delay_line_0.stop_strong.t5 a_9330_16954.t28 VGND.t137 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X530 VDPWR.t52 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 tdc_0.vernier_delay_line_0.start_pos.t3 VDPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X531 VGND.t118 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X532 VGND.t457 tdc_0.vernier_delay_line_0.stop_strong.t63 a_10958_25646.t9 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X533 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 VGND.t232 VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X534 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t274 VDPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X535 a_12420_35162# a_12310_35116# uo_out[5].t3 VDPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X536 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 uio_in[0].t4 VGND.t187 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X537 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 a_10108_37672.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X538 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.start_neg.t12 VDPWR.t66 VDPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X539 VGND.t458 tdc_0.vernier_delay_line_0.stop_strong.t64 a_10958_34774.t5 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X540 tdc_0.start_buffer_0.start_buff.t0 a_7140_10670# VGND.t147 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X541 VDPWR.t338 ui_in[6].t5 a_24240_18144# VDPWR.t337 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X542 tdc_0.vernier_delay_line_0.stop_strong.t21 a_9330_16954.t29 VDPWR.t150 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X543 VGND.t497 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VGND.t496 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X544 VDPWR.t189 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VDPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X545 VDPWR.t587 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 a_12310_25988# VDPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X546 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VDPWR.t508 VDPWR.t507 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X547 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 ui_in[4].t5 VGND.t223 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X548 VGND.t282 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X549 tdc_0.start_buffer_0.start_delay.t0 tdc_0.start_buffer_0.start_buff.t18 VGND.t379 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X550 VDPWR.t446 VDPWR.t444 a_15680_15464# VDPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X551 VGND.t284 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 a_25060_12248# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X552 a_15680_11634# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VDPWR.t373 VDPWR.t372 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X553 VDPWR.t238 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 a_12310_32834# VDPWR.t237 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X554 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X555 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_3.in.t5 a_24240_17262# VDPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X556 a_24240_11366# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VDPWR.t328 VDPWR.t327 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X557 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 VDPWR.t471 VDPWR.t470 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X558 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 VGND.t388 VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X559 a_23820_8460# input_stage_andpwr_0.fine_delay_unit_1.in VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X560 VGND.t415 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X561 variable_delay_short_0.in a_23820_8460# VDPWR.t223 VDPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X562 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VGND.t418 VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X563 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 VDPWR.t290 VDPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X564 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in.t5 a_24240_14314# VDPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X565 uo_out[0].t3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t346 VDPWR.t345 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X566 variable_delay_short_0.variable_delay_unit_1.in.t1 variable_delay_short_0.in VDPWR.t589 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X567 VGND.t82 tdc_0.vernier_delay_line_0.start_neg.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X568 variable_delay_dummy_0.out variable_delay_dummy_0.variable_delay_unit_1.in.t4 a_15680_11634# VDPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X569 a_10108_39954.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 a_10958_39338.t9 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X570 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward.t3 a_24240_26106# VDPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X571 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VDPWR.t441 VDPWR.t443 VDPWR.t442 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X572 variable_delay_dummy_0.in a_15322_8490# VGND.t83 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X573 uo_out[3].t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t183 VDPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X574 a_10958_25646.t8 tdc_0.vernier_delay_line_0.stop_strong.t65 VGND.t443 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X575 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 VGND.t177 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X576 input_stage_andpwr_0.fine_delay_unit_0.in input_stage_andpwr_0.nand_gate_0.out ua[0].t3 ua[0].t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X577 VGND.t471 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37444# VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X578 VGND.t511 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X579 VDPWR.t288 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 VDPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X580 a_10108_39954.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 a_10958_39338.t8 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X581 a_10958_37056.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 a_10108_37672.t2 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X582 a_12420_30598# a_12310_30552# uo_out[3].t3 VDPWR.t596 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X583 a_9330_14054# a_9330_13764# VDPWR.t81 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X584 a_13254_26412# uo_out[1].t5 VGND.t238 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X585 VDPWR.t380 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 VDPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X586 VGND.t317 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X587 a_9330_15504# a_9330_15214# VDPWR.t482 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X588 a_9330_16954.t5 a_9330_15794# VDPWR.t555 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X589 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 VDPWR.t40 VDPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X590 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t66 VDPWR.t489 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X591 tdc_0.vernier_delay_line_0.stop_strong.t20 a_9330_16954.t30 VDPWR.t403 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X592 a_25060_21092# variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X593 VGND.t499 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 a_12310_28270# VGND.t498 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X594 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 VDPWR.t234 VDPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X595 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 a_10108_28016# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X596 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 VDPWR.t330 VDPWR.t329 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X597 VGND.t441 tdc_0.vernier_delay_line_0.stop_strong.t67 a_10958_37056.t5 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X598 a_13254_32880# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 uo_out[4].t3 VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X599 a_10108_26262.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X600 ua[0].t4 VDPWR.t624 input_stage_andpwr_0.nand_gate_0.out ua[0].t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X601 tdc_0.vernier_delay_line_0.stop_strong.t19 a_9330_16954.t31 VDPWR.t404 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X602 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 VDPWR.t152 VDPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X603 VGND.t193 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 a_25060_24040# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X604 VGND.t347 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 a_12310_37398# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X605 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VGND.t263 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X606 variable_delay_short_0.variable_delay_unit_1.in.t0 variable_delay_short_0.in VGND.t548 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X607 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 VDPWR.t209 VDPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X608 VGND.t25 input_stage_andpwr_0.fine_delay_unit_1.in a_24790_8314# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X609 VGND.t349 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_23752# VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X610 a_12420_24130# uo_out[0].t5 VDPWR.t389 VDPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X611 VDPWR.t569 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 VDPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X612 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 a_10958_37056.t12 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X613 a_15322_7112# input_stage_0.fine_delay_unit_0.in a_16292_6702# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X614 VGND.t533 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_32880# VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X615 tdc_0.vernier_delay_line_0.stop_strong.t4 a_9330_16954.t32 VGND.t354 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X616 a_10958_34774.t4 tdc_0.vernier_delay_line_0.stop_strong.t68 VGND.t442 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X617 VGND.t320 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 a_16500_12516# VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X618 VDPWR.t158 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 VDPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X619 a_12420_33258# uo_out[4].t5 VDPWR.t522 VDPWR.t521 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X620 VDPWR.t394 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 VDPWR.t393 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X621 VGND.t412 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X622 uo_out[5].t2 a_12310_35116# VGND.t473 VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X623 a_10108_26262.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 a_10958_25646.t2 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X624 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 a_10108_33108.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X625 a_10958_27928.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 a_10108_28016# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X626 a_12420_40104# uo_out[7].t5 VDPWR.t218 VDPWR.t217 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X627 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 VDPWR.t284 VDPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X628 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VDPWR.t571 VDPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X629 a_13254_26034# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 uo_out[1].t2 VGND.t467 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X630 a_16292_6702# input_stage_0.fine_delay_unit_0.in a_15322_7112# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X631 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VDPWR.t583 VDPWR.t582 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X632 VGND.t357 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 a_25060_15196# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X633 a_10958_34774.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 a_10108_34862# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X634 variable_delay_dummy_0.variable_delay_unit_1.in.t1 variable_delay_dummy_0.in VDPWR.t485 VDPWR.t442 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X635 a_13254_35540# uo_out[5].t5 VGND.t257 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X636 VGND.t439 tdc_0.vernier_delay_line_0.stop_strong.t69 a_10958_32492.t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X637 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12308_31014# a_12420_30976# VDPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X638 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 VDPWR.t431 VDPWR.t430 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X639 a_10958_25646.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 a_10108_26262.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X640 input_stage_0.fine_delay_unit_1.in a_15322_7112# VGND.t416 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X641 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 VGND.t329 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X642 VGND.t216 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X643 VGND.t285 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 a_25060_12248# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X644 a_15680_11634# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VDPWR.t100 VDPWR.t99 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X645 a_10958_27928.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 a_10108_28016# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X646 a_10108_26262.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 a_10958_25646.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X647 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 VDPWR.t585 VDPWR.t584 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X648 VGND.t98 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 a_12310_23706# VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X649 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 VDPWR.t548 VDPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X650 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X651 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X652 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 a_10108_37144# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X653 VGND.t440 tdc_0.vernier_delay_line_0.stop_strong.t70 a_10958_30210.t1 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X654 VDPWR.t197 uio_in[0].t5 a_24240_12248# VDPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X655 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 tdc_0.start_buffer_0.start_buff.t19 VDPWR.t421 VDPWR.t420 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X656 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 VGND.t430 VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X657 VGND.t287 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 a_12310_30552# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X658 a_16500_12516# variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X659 a_10958_32492.t5 tdc_0.vernier_delay_line_0.stop_strong.t71 VGND.t436 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X660 VDPWR.t32 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12420_39726# VDPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X661 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 VGND.t293 VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X662 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 VDPWR.t76 VDPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X663 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 a_10958_23364.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X664 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.in.t4 a_25060_23158# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X665 a_16292_8344# input_stage_0.fine_delay_unit_1.in a_16292_8080# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X666 a_10958_39338.t4 tdc_0.vernier_delay_line_0.stop_strong.t72 VGND.t438 VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X667 a_24790_6672# input_stage_andpwr_0.fine_delay_unit_0.in a_23820_7082# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X668 VDPWR.t576 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X669 a_9330_14924# a_9330_14634# VGND.t549 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X670 VGND.t487 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X671 VDPWR.t366 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 VDPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X672 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t261 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X673 input_stage_0.nand_gate_0.out uio_in[5].t0 a_16786_5138# VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X674 VGND.t432 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X675 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_4.in.t4 a_25060_20210# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X676 a_10958_32492.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 a_10108_33108.t2 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X677 VDPWR.t213 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 VDPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X678 VGND.t243 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X679 VGND.t435 tdc_0.vernier_delay_line_0.stop_strong.t73 a_10958_30210.t0 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X680 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X681 a_9330_16954.t0 a_9330_15794# VGND.t525 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X682 VDPWR.t487 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 VDPWR.t486 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X683 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VDPWR.t46 VDPWR.t45 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X684 tdc_0.start_buffer_0.start_buff.t4 a_7140_10670# VDPWR.t159 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X685 VDPWR.t488 tdc_0.vernier_delay_line_0.stop_strong.t74 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X686 VGND.t378 tdc_0.start_buffer_0.start_buff.t20 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X687 VDPWR.t276 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 VDPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X688 tdc_0.vernier_delay_line_0.stop_strong.t3 a_9330_16954.t33 VGND.t134 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X689 tdc_0.start_buffer_0.start_delay.t4 tdc_0.start_buffer_0.start_buff.t21 VDPWR.t83 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X690 tdc_0.vernier_delay_line_0.stop_strong.t2 a_9330_16954.t34 VGND.t135 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X691 VGND.t38 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X692 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X693 VGND.t327 tdc_0.vernier_delay_line_0.stop_strong.t75 a_10958_23364.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X694 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 tdc_0.start_buffer_0.start_delay.t13 VDPWR.t201 VDPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X695 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 VGND.t515 VGND.t514 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X696 VGND.t104 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X697 a_13254_30976# uo_out[3].t5 VGND.t340 VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X698 tdc_0.vernier_delay_line_0.stop_strong.t18 a_9330_16954.t35 VDPWR.t147 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X699 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t76 VDPWR.t378 VDPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X700 VGND.t69 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X701 VGND.t519 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X702 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 VDPWR.t310 VDPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X703 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VGND.t175 VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X704 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 a_10108_23452# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X705 tdc_0.start_buffer_0.start_delay.t3 tdc_0.start_buffer_0.start_buff.t22 VGND.t376 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X706 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 VGND.t122 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X707 VGND.t428 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X708 a_10958_37056.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 a_10108_37144# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X709 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VGND.t168 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X710 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 a_10108_32580# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X711 VDPWR.t50 tdc_0.start_buffer_0.start_delay.t14 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 VDPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X712 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 VGND.t322 VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X713 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 VDPWR.t377 VDPWR.t376 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X714 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in.t4 a_25060_11366# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X715 a_24240_21092# variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out VDPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X716 VGND.t543 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 a_16500_15464# VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X717 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 VGND.t255 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X718 VDPWR.t478 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X719 VDPWR.t30 ui_in[4].t6 a_24240_24040# VDPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X720 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VGND.t61 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X721 VDPWR.t312 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 VDPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X722 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t347 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X723 VGND.t492 ui_in[1].t0 a_24790_6936# VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X724 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 a_10958_32492.t10 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X725 VDPWR.t119 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X726 a_16500_11634# VDPWR.t625 VGND.t398 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X727 VDPWR.t364 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VDPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X728 a_15322_7112# input_stage_0.fine_delay_unit_0.in VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X729 VDPWR.t538 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 VDPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X730 a_12420_28316# a_12310_28270# uo_out[2].t3 VDPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X731 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 a_10958_25646.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X732 VGND.t331 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X733 a_12420_37822# uo_out[6].t5 VDPWR.t494 VDPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X734 VDPWR.t107 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 VDPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X735 a_25060_14314# ui_in[7].t6 VGND.t123 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X736 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 tdc_0.start_buffer_0.start_delay.t15 VGND.t367 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X737 VGND.t324 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X738 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 VDPWR.t48 VDPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X739 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 a_10958_32492.t11 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X740 variable_delay_dummy_0.out variable_delay_dummy_0.variable_delay_unit_1.in.t5 a_16500_11634# VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X741 a_7140_10670# variable_delay_dummy_0.out VGND.t413 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X742 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X743 a_25060_11366# uio_in[0].t6 VGND.t362 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X744 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12308_28732# a_12420_28694# VDPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X745 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 VDPWR.t175 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X746 VDPWR.t578 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 a_12310_39680# VDPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X747 VDPWR.t259 tdc_0.vernier_delay_line_0.stop_strong.t77 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X748 VDPWR.t94 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 tdc_0.vernier_delay_line_0.start_neg.t5 VDPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X749 VDPWR.t211 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26034# VDPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X750 a_10958_23364.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 a_10108_23452# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X751 a_9330_14924# a_9330_14634# VDPWR.t594 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X752 VDPWR.t135 ui_in[7].t7 a_24240_15196# VDPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X753 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X754 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 VGND.t313 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X755 VGND.t236 tdc_0.vernier_delay_line_0.stop_strong.t78 a_10958_39338.t3 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X756 a_13254_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 uo_out[7].t1 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X757 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.start_pos.t14 VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X758 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out VGND.t295 VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X759 VDPWR.t440 VDPWR.t438 a_15680_12516# VDPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X760 a_9330_16954.t4 a_9330_15794# VDPWR.t554 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X761 a_10958_32492.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 a_10108_32580# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X762 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 VGND.t90 VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X763 VDPWR.t419 uio_in[0].t7 a_24240_12248# VDPWR.t418 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X764 VGND.t397 VDPWR.t626 a_25060_26106# VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X765 tdc_0.vernier_delay_line_0.stop_strong.t17 a_9330_16954.t36 VDPWR.t601 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X766 tdc_0.vernier_delay_line_0.stop_strong.t16 a_9330_16954.t37 VDPWR.t602 VDPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X767 tdc_0.vernier_delay_line_0.start_pos.t0 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 VGND.t173 VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X768 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X769 uo_out[7].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t498 VDPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X770 VDPWR.t44 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 VDPWR.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X771 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t144 VDPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X772 VGND.t34 ui_in[4].t7 a_25060_23158# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X773 VDPWR.t115 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VDPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X774 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 VDPWR.t253 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X775 VDPWR.t247 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X776 a_24240_26988# VDPWR.t435 VDPWR.t437 VDPWR.t436 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X777 a_10108_30826.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 a_10958_30210.t5 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X778 VGND.t517 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X779 tdc_0.vernier_delay_line_0.start_neg.t2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X780 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.in.t5 a_24240_23158# VDPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X781 VDPWR.t401 tdc_0.vernier_delay_line_0.stop_strong.t79 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X782 VDPWR.t177 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 VDPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X783 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t203 VDPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X784 VGND.t20 tdc_0.vernier_delay_line_0.start_pos.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X785 a_12420_37444# a_12310_37398# uo_out[6].t1 VDPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X786 VGND.t422 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X787 tdc_0.vernier_delay_line_0.stop_strong.t1 a_9330_16954.t38 VGND.t556 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X788 VGND.t375 tdc_0.start_buffer_0.start_buff.t23 tdc_0.start_buffer_0.start_delay.t2 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X789 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_4.in.t5 a_24240_20210# VDPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X790 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t146 VDPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X791 VGND.t185 ui_in[6].t6 a_25060_17262# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X792 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VDPWR.t298 VDPWR.t297 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X793 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t80 VDPWR.t402 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X794 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 VGND.t55 VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X795 VDPWR.t228 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VDPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X796 VDPWR.t249 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 a_12310_35116# VDPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X797 VGND.t495 uio_in[2].t0 a_16292_6966# VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X798 VGND.t445 tdc_0.vernier_delay_line_0.stop_strong.t81 a_10958_27928.t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X799 VGND.t67 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X800 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 VGND.t424 VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X801 VDPWR.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35162# VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X802 VDPWR.t268 tdc_0.vernier_delay_line_0.start_neg.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 VDPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X803 VGND.t536 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X804 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 VDPWR.t191 VDPWR.t190 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X805 uo_out[1].t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t205 VDPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X806 a_25060_17262# ui_in[6].t7 VGND.t186 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X807 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 VGND.t165 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X808 a_15680_15464# VDPWR.t432 VDPWR.t434 VDPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X809 a_10958_37056.t4 tdc_0.vernier_delay_line_0.stop_strong.t82 VGND.t446 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X810 VDPWR.t396 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 VDPWR.t395 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X811 a_16500_14582# VDPWR.t627 VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X812 VGND.t273 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X813 uo_out[4].t2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t357 VDPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X814 a_10958_27928.t5 tdc_0.vernier_delay_line_0.stop_strong.t83 VGND.t144 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X815 uo_out[2].t2 a_12310_28270# VGND.t551 VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X816 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in.t5 a_24240_11366# VDPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X817 VGND.t386 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X818 VGND.t145 tdc_0.vernier_delay_line_0.stop_strong.t84 a_10958_27928.t4 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X819 a_16500_11634# VDPWR.t628 VGND.t393 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X820 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VGND.t212 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X821 a_12420_23752# a_12310_23706# uo_out[0].t1 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X822 VDPWR.t86 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 VDPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X823 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.start_neg.t15 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X824 VGND.t444 tdc_0.vernier_delay_line_0.stop_strong.t85 a_10958_25646.t7 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X825 a_9330_15794# a_9330_15504# VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X826 VGND.t353 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X827 a_13254_28694# uo_out[2].t5 VGND.t96 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X828 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X829 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t86 VDPWR.t490 VDPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X830 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12308_24168# a_12420_24130# VDPWR.t468 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X831 input_stage_andpwr_0.fine_delay_unit_1.in a_23820_7082# VDPWR.t179 VDPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X832 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 VGND.t220 VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X833 VDPWR.t534 uio_in[5].t1 input_stage_0.nand_gate_0.out VDPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X834 VDPWR.t154 tdc_0.vernier_delay_line_0.stop_strong.t87 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X835 tdc_0.vernier_delay_line_0.stop_strong.t0 a_9330_16954.t39 VGND.t280 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 552.84
R1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 552.84
R2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 552.84
R3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 552.84
R4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 539.841
R5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 539.841
R6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 539.841
R7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 539.841
R8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 215.293
R9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 215.293
R10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 215.293
R11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 215.293
R12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 166.468
R13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 166.149
R14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 165.8
R15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 165.8
R16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 85.1574
R17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 83.8097
R18 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 83.8097
R19 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 83.7172
R20 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 74.288
R21 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 67.7574
R22 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 36.1505
R23 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 36.1505
R24 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 34.5438
R25 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 34.5438
R26 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 17.4005
R27 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 17.4005
R28 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 16.09
R29 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 11.8364
R30 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 9.52217
R31 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 9.52217
R32 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 5.96628
R33 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 5.83219
R34 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 5.74235
R35 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 5.49235
R36 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 1.44072
R37 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 1.32081
R38 VDPWR.n1186 VDPWR.n1185 2207.5
R39 VDPWR.n1202 VDPWR.n1201 2207.5
R40 VDPWR.n1218 VDPWR.n1217 2207.5
R41 VDPWR.n1234 VDPWR.n1233 2207.5
R42 VDPWR.n1250 VDPWR.n1249 2207.5
R43 VDPWR.n1266 VDPWR.n1265 2207.5
R44 VDPWR.n1282 VDPWR.n1281 2207.5
R45 VDPWR.n1298 VDPWR.n1297 2207.5
R46 VDPWR.n1376 VDPWR.n1350 2207.5
R47 VDPWR.n1396 VDPWR.n1350 2207.5
R48 VDPWR.n1398 VDPWR.n1349 2207.5
R49 VDPWR.n1404 VDPWR.n1349 2207.5
R50 VDPWR.n1402 VDPWR.n1334 2207.5
R51 VDPWR.n1424 VDPWR.n1334 2207.5
R52 VDPWR.n1426 VDPWR.n1333 2207.5
R53 VDPWR.n1432 VDPWR.n1333 2207.5
R54 VDPWR.n1430 VDPWR.n1318 2207.5
R55 VDPWR.n1452 VDPWR.n1318 2207.5
R56 VDPWR.n1454 VDPWR.n1317 2207.5
R57 VDPWR.n983 VDPWR.n977 2106.47
R58 VDPWR.n1001 VDPWR.n995 2106.47
R59 VDPWR.n1019 VDPWR.n1013 2106.47
R60 VDPWR.n1037 VDPWR.n1031 2106.47
R61 VDPWR.n1055 VDPWR.n1049 2106.47
R62 VDPWR.n1073 VDPWR.n1067 2106.47
R63 VDPWR.n1091 VDPWR.n1085 2106.47
R64 VDPWR.n1109 VDPWR.n1103 2106.47
R65 VDPWR.n979 VDPWR.n978 2101.76
R66 VDPWR.n997 VDPWR.n996 2101.76
R67 VDPWR.n1015 VDPWR.n1014 2101.76
R68 VDPWR.n1033 VDPWR.n1032 2101.76
R69 VDPWR.n1051 VDPWR.n1050 2101.76
R70 VDPWR.n1069 VDPWR.n1068 2101.76
R71 VDPWR.n1087 VDPWR.n1086 2101.76
R72 VDPWR.n1105 VDPWR.n1104 2101.76
R73 VDPWR.n1170 VDPWR.n1165 2093.75
R74 VDPWR.n1371 VDPWR.n1365 2093.75
R75 VDPWR.n1175 VDPWR.n1166 2088.75
R76 VDPWR.n1380 VDPWR.n1366 2088.75
R77 VDPWR.n1187 VDPWR.n1185 2070
R78 VDPWR.n1203 VDPWR.n1201 2070
R79 VDPWR.n1219 VDPWR.n1217 2070
R80 VDPWR.n1235 VDPWR.n1233 2070
R81 VDPWR.n1251 VDPWR.n1249 2070
R82 VDPWR.n1267 VDPWR.n1265 2070
R83 VDPWR.n1283 VDPWR.n1281 2070
R84 VDPWR.n1299 VDPWR.n1297 2070
R85 VDPWR.n1456 VDPWR.n1317 2070
R86 VDPWR.n201 VDPWR.n198 1689.71
R87 VDPWR.n467 VDPWR.n198 1689.71
R88 VDPWR.n471 VDPWR.n197 1689.71
R89 VDPWR.n471 VDPWR.n196 1689.71
R90 VDPWR.n225 VDPWR.n222 1689.71
R91 VDPWR.n441 VDPWR.n222 1689.71
R92 VDPWR.n445 VDPWR.n221 1689.71
R93 VDPWR.n445 VDPWR.n220 1689.71
R94 VDPWR.n249 VDPWR.n246 1689.71
R95 VDPWR.n415 VDPWR.n246 1689.71
R96 VDPWR.n419 VDPWR.n245 1689.71
R97 VDPWR.n419 VDPWR.n244 1689.71
R98 VDPWR.n273 VDPWR.n270 1689.71
R99 VDPWR.n389 VDPWR.n270 1689.71
R100 VDPWR.n393 VDPWR.n269 1689.71
R101 VDPWR.n393 VDPWR.n268 1689.71
R102 VDPWR.n297 VDPWR.n294 1689.71
R103 VDPWR.n363 VDPWR.n294 1689.71
R104 VDPWR.n367 VDPWR.n293 1689.71
R105 VDPWR.n367 VDPWR.n292 1689.71
R106 VDPWR.n321 VDPWR.n318 1689.71
R107 VDPWR.n329 VDPWR.n318 1689.71
R108 VDPWR.n333 VDPWR.n317 1689.71
R109 VDPWR.n333 VDPWR.n316 1689.71
R110 VDPWR.n32 VDPWR.n29 1689.71
R111 VDPWR.n98 VDPWR.n29 1689.71
R112 VDPWR.n102 VDPWR.n28 1689.71
R113 VDPWR.n102 VDPWR.n27 1689.71
R114 VDPWR.n56 VDPWR.n53 1689.71
R115 VDPWR.n64 VDPWR.n53 1689.71
R116 VDPWR.n68 VDPWR.n52 1689.71
R117 VDPWR.n68 VDPWR.n51 1689.71
R118 VDPWR.n683 VDPWR.n516 1508.99
R119 VDPWR.n666 VDPWR.n521 1508.99
R120 VDPWR.n649 VDPWR.n526 1508.99
R121 VDPWR.n632 VDPWR.n531 1508.99
R122 VDPWR.n615 VDPWR.n536 1508.99
R123 VDPWR.n598 VDPWR.n541 1508.99
R124 VDPWR.n581 VDPWR.n546 1508.99
R125 VDPWR.n564 VDPWR.n551 1508.99
R126 VDPWR.n980 VDPWR.n978 1450
R127 VDPWR.n998 VDPWR.n996 1450
R128 VDPWR.n1016 VDPWR.n1014 1450
R129 VDPWR.n1034 VDPWR.n1032 1450
R130 VDPWR.n1052 VDPWR.n1050 1450
R131 VDPWR.n1070 VDPWR.n1068 1450
R132 VDPWR.n1088 VDPWR.n1086 1450
R133 VDPWR.n1106 VDPWR.n1104 1450
R134 VDPWR.n1549 VDPWR.n164 1348.04
R135 VDPWR.n1171 VDPWR.n1165 1326.32
R136 VDPWR.n1372 VDPWR.n1365 1326.32
R137 VDPWR.n679 VDPWR.n677 1313.33
R138 VDPWR.n662 VDPWR.n660 1313.33
R139 VDPWR.n645 VDPWR.n643 1313.33
R140 VDPWR.n628 VDPWR.n626 1313.33
R141 VDPWR.n611 VDPWR.n609 1313.33
R142 VDPWR.n594 VDPWR.n592 1313.33
R143 VDPWR.n577 VDPWR.n575 1313.33
R144 VDPWR.n560 VDPWR.n558 1313.33
R145 VDPWR.n1489 VDPWR.n1468 1307.92
R146 VDPWR.n1507 VDPWR.n1500 1307.92
R147 VDPWR.n783 VDPWR.n689 1307.92
R148 VDPWR.n840 VDPWR.n782 1307.92
R149 VDPWR.n481 VDPWR.n187 1307.92
R150 VDPWR.n481 VDPWR.n188 1307.92
R151 VDPWR.n483 VDPWR.n185 1307.92
R152 VDPWR.n483 VDPWR.n184 1307.92
R153 VDPWR.n455 VDPWR.n211 1307.92
R154 VDPWR.n455 VDPWR.n212 1307.92
R155 VDPWR.n457 VDPWR.n209 1307.92
R156 VDPWR.n457 VDPWR.n208 1307.92
R157 VDPWR.n429 VDPWR.n235 1307.92
R158 VDPWR.n429 VDPWR.n236 1307.92
R159 VDPWR.n431 VDPWR.n233 1307.92
R160 VDPWR.n431 VDPWR.n232 1307.92
R161 VDPWR.n403 VDPWR.n259 1307.92
R162 VDPWR.n403 VDPWR.n260 1307.92
R163 VDPWR.n405 VDPWR.n257 1307.92
R164 VDPWR.n405 VDPWR.n256 1307.92
R165 VDPWR.n377 VDPWR.n283 1307.92
R166 VDPWR.n377 VDPWR.n284 1307.92
R167 VDPWR.n379 VDPWR.n281 1307.92
R168 VDPWR.n379 VDPWR.n280 1307.92
R169 VDPWR.n343 VDPWR.n307 1307.92
R170 VDPWR.n343 VDPWR.n308 1307.92
R171 VDPWR.n345 VDPWR.n305 1307.92
R172 VDPWR.n345 VDPWR.n304 1307.92
R173 VDPWR.n154 VDPWR.n153 1307.92
R174 VDPWR.n112 VDPWR.n18 1307.92
R175 VDPWR.n112 VDPWR.n19 1307.92
R176 VDPWR.n114 VDPWR.n16 1307.92
R177 VDPWR.n114 VDPWR.n15 1307.92
R178 VDPWR.n80 VDPWR.n39 1307.92
R179 VDPWR.n80 VDPWR.n40 1307.92
R180 VDPWR.n78 VDPWR.n42 1307.92
R181 VDPWR.n78 VDPWR.n43 1307.92
R182 VDPWR.n492 VDPWR.n178 1271.17
R183 VDPWR.n503 VDPWR.n172 1271.17
R184 VDPWR.n131 VDPWR.n9 1271.17
R185 VDPWR.n142 VDPWR.n3 1271.17
R186 VDPWR.n1517 VDPWR.n1488 1126.67
R187 VDPWR.n1491 VDPWR.n1490 1126.67
R188 VDPWR.n1493 VDPWR.n1492 1126.67
R189 VDPWR.n1495 VDPWR.n1494 1126.67
R190 VDPWR.n1497 VDPWR.n1496 1126.67
R191 VDPWR.n1499 VDPWR.n1498 1126.67
R192 VDPWR.n1515 VDPWR.n1502 1126.67
R193 VDPWR.n785 VDPWR.n784 1126.67
R194 VDPWR.n787 VDPWR.n786 1126.67
R195 VDPWR.n789 VDPWR.n788 1126.67
R196 VDPWR.n791 VDPWR.n790 1126.67
R197 VDPWR.n793 VDPWR.n792 1126.67
R198 VDPWR.n795 VDPWR.n794 1126.67
R199 VDPWR.n797 VDPWR.n796 1126.67
R200 VDPWR.n799 VDPWR.n798 1126.67
R201 VDPWR.n801 VDPWR.n800 1126.67
R202 VDPWR.n803 VDPWR.n802 1126.67
R203 VDPWR.n805 VDPWR.n804 1126.67
R204 VDPWR.n807 VDPWR.n806 1126.67
R205 VDPWR.n809 VDPWR.n808 1126.67
R206 VDPWR.n811 VDPWR.n810 1126.67
R207 VDPWR.n813 VDPWR.n812 1126.67
R208 VDPWR.n815 VDPWR.n814 1126.67
R209 VDPWR.n817 VDPWR.n816 1126.67
R210 VDPWR.n819 VDPWR.n818 1126.67
R211 VDPWR.n821 VDPWR.n820 1126.67
R212 VDPWR.n823 VDPWR.n822 1126.67
R213 VDPWR.n825 VDPWR.n824 1126.67
R214 VDPWR.n827 VDPWR.n826 1126.67
R215 VDPWR.n829 VDPWR.n828 1126.67
R216 VDPWR.n831 VDPWR.n830 1126.67
R217 VDPWR.n833 VDPWR.n832 1126.67
R218 VDPWR.n838 VDPWR.n837 1126.67
R219 VDPWR.n835 VDPWR.n834 1126.67
R220 VDPWR.n351 VDPWR.t456 628.097
R221 VDPWR.n120 VDPWR.t450 628.097
R222 VDPWR.n86 VDPWR.t459 628.097
R223 VDPWR.n352 VDPWR.t447 622.766
R224 VDPWR.n121 VDPWR.t438 622.766
R225 VDPWR.n87 VDPWR.t444 622.766
R226 VDPWR.n167 VDPWR.t624 564.04
R227 VDPWR.n156 VDPWR.n153 551.179
R228 VDPWR.n350 VDPWR.t465 543.053
R229 VDPWR.n119 VDPWR.t441 543.053
R230 VDPWR.n85 VDPWR.t453 543.053
R231 VDPWR.n351 VDPWR.t435 523.774
R232 VDPWR.n120 VDPWR.t462 523.774
R233 VDPWR.n86 VDPWR.t432 523.774
R234 VDPWR.n167 VDPWR.t621 511.623
R235 VDPWR.n1547 VDPWR.n164 485.663
R236 VDPWR.n482 VDPWR.n186 460.678
R237 VDPWR.n456 VDPWR.n210 460.678
R238 VDPWR.n430 VDPWR.n234 460.678
R239 VDPWR.n404 VDPWR.n258 460.678
R240 VDPWR.n378 VDPWR.n282 460.678
R241 VDPWR.n344 VDPWR.n306 460.678
R242 VDPWR.n113 VDPWR.n17 460.678
R243 VDPWR.n79 VDPWR.n41 460.678
R244 VDPWR.n180 VDPWR.n178 408.981
R245 VDPWR.n174 VDPWR.n172 408.981
R246 VDPWR.n11 VDPWR.n9 408.981
R247 VDPWR.n5 VDPWR.n3 408.981
R248 VDPWR.n682 VDPWR.n675 358.526
R249 VDPWR.n665 VDPWR.n658 358.526
R250 VDPWR.n648 VDPWR.n641 358.526
R251 VDPWR.n631 VDPWR.n624 358.526
R252 VDPWR.n614 VDPWR.n607 358.526
R253 VDPWR.n597 VDPWR.n590 358.526
R254 VDPWR.n580 VDPWR.n573 358.526
R255 VDPWR.n563 VDPWR.n556 358.526
R256 VDPWR.n469 VDPWR.n468 332.803
R257 VDPWR.n443 VDPWR.n442 332.803
R258 VDPWR.n417 VDPWR.n416 332.803
R259 VDPWR.n391 VDPWR.n390 332.803
R260 VDPWR.n365 VDPWR.n364 332.803
R261 VDPWR.n331 VDPWR.n330 332.803
R262 VDPWR.n100 VDPWR.n99 332.803
R263 VDPWR.n66 VDPWR.n65 332.803
R264 VDPWR.n495 VDPWR.n494 313.632
R265 VDPWR.n134 VDPWR.n133 313.632
R266 VDPWR.n506 VDPWR.n505 312.635
R267 VDPWR.n145 VDPWR.n144 312.635
R268 VDPWR.n353 VDPWR.t617 304.647
R269 VDPWR.n353 VDPWR.t623 304.647
R270 VDPWR.n122 VDPWR.t625 304.647
R271 VDPWR.n122 VDPWR.t628 304.647
R272 VDPWR.n88 VDPWR.t619 304.647
R273 VDPWR.n88 VDPWR.t627 304.647
R274 VDPWR.n674 VDPWR.n672 254.195
R275 VDPWR.n657 VDPWR.n655 254.195
R276 VDPWR.n640 VDPWR.n638 254.195
R277 VDPWR.n623 VDPWR.n621 254.195
R278 VDPWR.n606 VDPWR.n604 254.195
R279 VDPWR.n589 VDPWR.n587 254.195
R280 VDPWR.n572 VDPWR.n570 254.195
R281 VDPWR.n555 VDPWR.n553 254.195
R282 VDPWR.n1192 VDPWR.n1184 235.468
R283 VDPWR.n1208 VDPWR.n1200 235.468
R284 VDPWR.n1224 VDPWR.n1216 235.468
R285 VDPWR.n1240 VDPWR.n1232 235.468
R286 VDPWR.n1256 VDPWR.n1248 235.468
R287 VDPWR.n1272 VDPWR.n1264 235.468
R288 VDPWR.n1288 VDPWR.n1280 235.468
R289 VDPWR.n1304 VDPWR.n1296 235.468
R290 VDPWR.n1394 VDPWR.n1355 235.468
R291 VDPWR.n1395 VDPWR.n1394 235.468
R292 VDPWR.n1409 VDPWR.n1348 235.468
R293 VDPWR.n1409 VDPWR.n1343 235.468
R294 VDPWR.n1422 VDPWR.n1339 235.468
R295 VDPWR.n1423 VDPWR.n1422 235.468
R296 VDPWR.n1437 VDPWR.n1332 235.468
R297 VDPWR.n1437 VDPWR.n1327 235.468
R298 VDPWR.n1450 VDPWR.n1323 235.468
R299 VDPWR.n1451 VDPWR.n1450 235.468
R300 VDPWR.n1461 VDPWR.n1316 235.468
R301 VDPWR.n985 VDPWR.n976 224.69
R302 VDPWR.n1003 VDPWR.n994 224.69
R303 VDPWR.n1021 VDPWR.n1012 224.69
R304 VDPWR.n1039 VDPWR.n1030 224.69
R305 VDPWR.n1057 VDPWR.n1048 224.69
R306 VDPWR.n1075 VDPWR.n1066 224.69
R307 VDPWR.n1093 VDPWR.n1084 224.69
R308 VDPWR.n1111 VDPWR.n1102 224.69
R309 VDPWR.n984 VDPWR.n970 224.189
R310 VDPWR.n1002 VDPWR.n966 224.189
R311 VDPWR.n1020 VDPWR.n962 224.189
R312 VDPWR.n1038 VDPWR.n958 224.189
R313 VDPWR.n1056 VDPWR.n954 224.189
R314 VDPWR.n1074 VDPWR.n950 224.189
R315 VDPWR.n1092 VDPWR.n946 224.189
R316 VDPWR.n1110 VDPWR.n942 224.189
R317 VDPWR.n1169 VDPWR.n1164 223.333
R318 VDPWR.n1370 VDPWR.n1364 223.333
R319 VDPWR.n1176 VDPWR.n1159 222.8
R320 VDPWR.n1381 VDPWR.n1359 222.8
R321 VDPWR.n350 VDPWR.t615 221.72
R322 VDPWR.n119 VDPWR.t620 221.72
R323 VDPWR.n85 VDPWR.t616 221.72
R324 VDPWR.n1192 VDPWR.n1154 220.8
R325 VDPWR.n1208 VDPWR.n1149 220.8
R326 VDPWR.n1224 VDPWR.n1144 220.8
R327 VDPWR.n1240 VDPWR.n1139 220.8
R328 VDPWR.n1256 VDPWR.n1134 220.8
R329 VDPWR.n1272 VDPWR.n1129 220.8
R330 VDPWR.n1288 VDPWR.n1124 220.8
R331 VDPWR.n1304 VDPWR.n1119 220.8
R332 VDPWR.n1461 VDPWR.n1311 220.8
R333 VDPWR.n125 VDPWR.n119 219.549
R334 VDPWR.n91 VDPWR.n85 219.531
R335 VDPWR.n356 VDPWR.n350 219.526
R336 VDPWR.n353 VDPWR.t626 202.44
R337 VDPWR.n122 VDPWR.t622 202.44
R338 VDPWR.n88 VDPWR.t618 202.44
R339 VDPWR.n681 VDPWR.n680 185.162
R340 VDPWR.n664 VDPWR.n663 185.162
R341 VDPWR.n647 VDPWR.n646 185.162
R342 VDPWR.n630 VDPWR.n629 185.162
R343 VDPWR.n613 VDPWR.n612 185.162
R344 VDPWR.n596 VDPWR.n595 185.162
R345 VDPWR.n579 VDPWR.n578 185.162
R346 VDPWR.n562 VDPWR.n561 185.162
R347 VDPWR.n682 VDPWR.n681 185
R348 VDPWR.n665 VDPWR.n664 185
R349 VDPWR.n648 VDPWR.n647 185
R350 VDPWR.n631 VDPWR.n630 185
R351 VDPWR.n614 VDPWR.n613 185
R352 VDPWR.n597 VDPWR.n596 185
R353 VDPWR.n580 VDPWR.n579 185
R354 VDPWR.n563 VDPWR.n562 185
R355 VDPWR.n1490 VDPWR.n1468 181.25
R356 VDPWR.n1490 VDPWR.n1470 181.25
R357 VDPWR.n1492 VDPWR.n1470 181.25
R358 VDPWR.n1492 VDPWR.n1475 181.25
R359 VDPWR.n1494 VDPWR.n1475 181.25
R360 VDPWR.n1494 VDPWR.n1477 181.25
R361 VDPWR.n1496 VDPWR.n1477 181.25
R362 VDPWR.n1496 VDPWR.n1482 181.25
R363 VDPWR.n1498 VDPWR.n1482 181.25
R364 VDPWR.n1498 VDPWR.n1484 181.25
R365 VDPWR.n1488 VDPWR.n1484 181.25
R366 VDPWR.n1505 VDPWR.n1488 181.25
R367 VDPWR.n1505 VDPWR.n1502 181.25
R368 VDPWR.n1507 VDPWR.n1502 181.25
R369 VDPWR.n784 VDPWR.n689 181.25
R370 VDPWR.n784 VDPWR.n691 181.25
R371 VDPWR.n786 VDPWR.n691 181.25
R372 VDPWR.n786 VDPWR.n696 181.25
R373 VDPWR.n788 VDPWR.n696 181.25
R374 VDPWR.n788 VDPWR.n698 181.25
R375 VDPWR.n790 VDPWR.n698 181.25
R376 VDPWR.n790 VDPWR.n703 181.25
R377 VDPWR.n792 VDPWR.n703 181.25
R378 VDPWR.n792 VDPWR.n705 181.25
R379 VDPWR.n794 VDPWR.n705 181.25
R380 VDPWR.n794 VDPWR.n710 181.25
R381 VDPWR.n796 VDPWR.n710 181.25
R382 VDPWR.n796 VDPWR.n712 181.25
R383 VDPWR.n798 VDPWR.n712 181.25
R384 VDPWR.n798 VDPWR.n717 181.25
R385 VDPWR.n800 VDPWR.n717 181.25
R386 VDPWR.n800 VDPWR.n719 181.25
R387 VDPWR.n802 VDPWR.n719 181.25
R388 VDPWR.n802 VDPWR.n724 181.25
R389 VDPWR.n804 VDPWR.n724 181.25
R390 VDPWR.n804 VDPWR.n726 181.25
R391 VDPWR.n806 VDPWR.n726 181.25
R392 VDPWR.n806 VDPWR.n731 181.25
R393 VDPWR.n808 VDPWR.n731 181.25
R394 VDPWR.n808 VDPWR.n733 181.25
R395 VDPWR.n810 VDPWR.n733 181.25
R396 VDPWR.n810 VDPWR.n738 181.25
R397 VDPWR.n812 VDPWR.n738 181.25
R398 VDPWR.n812 VDPWR.n740 181.25
R399 VDPWR.n814 VDPWR.n740 181.25
R400 VDPWR.n814 VDPWR.n745 181.25
R401 VDPWR.n816 VDPWR.n745 181.25
R402 VDPWR.n816 VDPWR.n747 181.25
R403 VDPWR.n818 VDPWR.n747 181.25
R404 VDPWR.n818 VDPWR.n752 181.25
R405 VDPWR.n820 VDPWR.n752 181.25
R406 VDPWR.n820 VDPWR.n754 181.25
R407 VDPWR.n822 VDPWR.n754 181.25
R408 VDPWR.n822 VDPWR.n759 181.25
R409 VDPWR.n824 VDPWR.n759 181.25
R410 VDPWR.n824 VDPWR.n761 181.25
R411 VDPWR.n826 VDPWR.n761 181.25
R412 VDPWR.n826 VDPWR.n766 181.25
R413 VDPWR.n828 VDPWR.n766 181.25
R414 VDPWR.n828 VDPWR.n768 181.25
R415 VDPWR.n830 VDPWR.n768 181.25
R416 VDPWR.n830 VDPWR.n773 181.25
R417 VDPWR.n832 VDPWR.n773 181.25
R418 VDPWR.n832 VDPWR.n775 181.25
R419 VDPWR.n837 VDPWR.n775 181.25
R420 VDPWR.n837 VDPWR.n780 181.25
R421 VDPWR.n834 VDPWR.n780 181.25
R422 VDPWR.n834 VDPWR.n782 181.25
R423 VDPWR.n465 VDPWR.n202 180.236
R424 VDPWR.n466 VDPWR.n465 180.236
R425 VDPWR.n472 VDPWR.n195 180.236
R426 VDPWR.n472 VDPWR.n191 180.236
R427 VDPWR.n439 VDPWR.n226 180.236
R428 VDPWR.n440 VDPWR.n439 180.236
R429 VDPWR.n446 VDPWR.n219 180.236
R430 VDPWR.n446 VDPWR.n215 180.236
R431 VDPWR.n413 VDPWR.n250 180.236
R432 VDPWR.n414 VDPWR.n413 180.236
R433 VDPWR.n420 VDPWR.n243 180.236
R434 VDPWR.n420 VDPWR.n239 180.236
R435 VDPWR.n387 VDPWR.n274 180.236
R436 VDPWR.n388 VDPWR.n387 180.236
R437 VDPWR.n394 VDPWR.n267 180.236
R438 VDPWR.n394 VDPWR.n263 180.236
R439 VDPWR.n361 VDPWR.n298 180.236
R440 VDPWR.n362 VDPWR.n361 180.236
R441 VDPWR.n368 VDPWR.n291 180.236
R442 VDPWR.n368 VDPWR.n287 180.236
R443 VDPWR.n327 VDPWR.n322 180.236
R444 VDPWR.n328 VDPWR.n327 180.236
R445 VDPWR.n334 VDPWR.n315 180.236
R446 VDPWR.n334 VDPWR.n311 180.236
R447 VDPWR.n96 VDPWR.n33 180.236
R448 VDPWR.n97 VDPWR.n96 180.236
R449 VDPWR.n103 VDPWR.n26 180.236
R450 VDPWR.n103 VDPWR.n22 180.236
R451 VDPWR.n62 VDPWR.n57 180.236
R452 VDPWR.n63 VDPWR.n62 180.236
R453 VDPWR.n69 VDPWR.n50 180.236
R454 VDPWR.n69 VDPWR.n46 180.236
R455 VDPWR.n1191 VDPWR.n1190 171.775
R456 VDPWR.n1207 VDPWR.n1206 171.775
R457 VDPWR.n1223 VDPWR.n1222 171.775
R458 VDPWR.n1239 VDPWR.n1238 171.775
R459 VDPWR.n1255 VDPWR.n1254 171.775
R460 VDPWR.n1271 VDPWR.n1270 171.775
R461 VDPWR.n1287 VDPWR.n1286 171.775
R462 VDPWR.n1303 VDPWR.n1302 171.775
R463 VDPWR.n1375 VDPWR.n1356 171.775
R464 VDPWR.n1408 VDPWR.n1407 171.775
R465 VDPWR.n1401 VDPWR.n1340 171.775
R466 VDPWR.n1436 VDPWR.n1435 171.775
R467 VDPWR.n1429 VDPWR.n1324 171.775
R468 VDPWR.n1460 VDPWR.n1459 171.775
R469 VDPWR.t384 VDPWR.n977 169.983
R470 VDPWR.t63 VDPWR.n995 169.983
R471 VDPWR.t397 VDPWR.n1013 169.983
R472 VDPWR.t145 VDPWR.n1031 169.983
R473 VDPWR.t184 VDPWR.n1049 169.983
R474 VDPWR.t319 VDPWR.n1067 169.983
R475 VDPWR.t202 VDPWR.n1085 169.983
R476 VDPWR.t273 VDPWR.n1103 169.983
R477 VDPWR VDPWR.n353 169.071
R478 VDPWR VDPWR.n122 169.071
R479 VDPWR VDPWR.n88 169.071
R480 VDPWR VDPWR.n352 166.244
R481 VDPWR VDPWR.n121 166.244
R482 VDPWR VDPWR.n87 166.244
R483 VDPWR.t577 VDPWR.n979 164.046
R484 VDPWR.t167 VDPWR.n997 164.046
R485 VDPWR.t248 VDPWR.n1015 164.046
R486 VDPWR.t237 VDPWR.n1033 164.046
R487 VDPWR.t155 VDPWR.n1051 164.046
R488 VDPWR.t324 VDPWR.n1069 164.046
R489 VDPWR.t586 VDPWR.n1087 164.046
R490 VDPWR.t599 VDPWR.n1105 164.046
R491 VDPWR.n201 VDPWR.t196 163.724
R492 VDPWR.t559 VDPWR.n197 163.724
R493 VDPWR.n225 VDPWR.t163 163.724
R494 VDPWR.t426 VDPWR.n221 163.724
R495 VDPWR.n249 VDPWR.t592 163.724
R496 VDPWR.t283 VDPWR.n245 163.724
R497 VDPWR.n273 VDPWR.t301 163.724
R498 VDPWR.t333 VDPWR.n269 163.724
R499 VDPWR.n297 VDPWR.t610 163.724
R500 VDPWR.t208 VDPWR.n293 163.724
R501 VDPWR.n321 VDPWR.t457 163.724
R502 VDPWR.t329 VDPWR.n317 163.724
R503 VDPWR.n32 VDPWR.t451 163.724
R504 VDPWR.t99 VDPWR.n28 163.724
R505 VDPWR.n56 VDPWR.t460 163.724
R506 VDPWR.t582 VDPWR.n52 163.724
R507 VDPWR.n168 VDPWR.n167 161.3
R508 VDPWR.n566 VDPWR.n565 160.959
R509 VDPWR.n583 VDPWR.n582 160.959
R510 VDPWR.n600 VDPWR.n599 160.959
R511 VDPWR.n617 VDPWR.n616 160.959
R512 VDPWR.n634 VDPWR.n633 160.959
R513 VDPWR.n651 VDPWR.n650 160.959
R514 VDPWR.n668 VDPWR.n667 160.959
R515 VDPWR.n685 VDPWR.n684 160.959
R516 VDPWR.n1171 VDPWR.n1164 158.292
R517 VDPWR.n1372 VDPWR.n1364 158.292
R518 VDPWR.n984 VDPWR.n972 154.667
R519 VDPWR.n1002 VDPWR.n968 154.667
R520 VDPWR.n1020 VDPWR.n964 154.667
R521 VDPWR.n1038 VDPWR.n960 154.667
R522 VDPWR.n1056 VDPWR.n956 154.667
R523 VDPWR.n1074 VDPWR.n952 154.667
R524 VDPWR.n1092 VDPWR.n948 154.667
R525 VDPWR.n1110 VDPWR.n944 154.667
R526 VDPWR.n680 VDPWR.n679 153.304
R527 VDPWR.n663 VDPWR.n662 153.304
R528 VDPWR.n646 VDPWR.n645 153.304
R529 VDPWR.n629 VDPWR.n628 153.304
R530 VDPWR.n612 VDPWR.n611 153.304
R531 VDPWR.n595 VDPWR.n594 153.304
R532 VDPWR.n578 VDPWR.n577 153.304
R533 VDPWR.n561 VDPWR.n560 153.304
R534 VDPWR.t470 VDPWR.n1170 151.868
R535 VDPWR.t547 VDPWR.n1186 151.868
R536 VDPWR.t194 VDPWR.n1202 151.868
R537 VDPWR.t61 VDPWR.n1218 151.868
R538 VDPWR.t281 VDPWR.n1234 151.868
R539 VDPWR.t293 VDPWR.n1250 151.868
R540 VDPWR.t526 VDPWR.n1266 151.868
R541 VDPWR.t108 VDPWR.n1282 151.868
R542 VDPWR.t12 VDPWR.n1298 151.868
R543 VDPWR.t14 VDPWR.n1371 151.868
R544 VDPWR.n1516 VDPWR.n1501 151.03
R545 VDPWR.n468 VDPWR.t199 145.224
R546 VDPWR.t606 VDPWR.n469 145.224
R547 VDPWR.n442 VDPWR.t509 145.224
R548 VDPWR.t491 VDPWR.n443 145.224
R549 VDPWR.n416 VDPWR.t558 145.224
R550 VDPWR.t171 VDPWR.n417 145.224
R551 VDPWR.n390 VDPWR.t226 145.224
R552 VDPWR.t129 VDPWR.n391 145.224
R553 VDPWR.n364 VDPWR.t3 145.224
R554 VDPWR.t390 VDPWR.n365 145.224
R555 VDPWR.n330 VDPWR.t112 145.224
R556 VDPWR.t520 VDPWR.n331 145.224
R557 VDPWR.n99 VDPWR.t511 145.224
R558 VDPWR.t102 VDPWR.n100 145.224
R559 VDPWR.n65 VDPWR.t113 145.224
R560 VDPWR.t138 VDPWR.n66 145.224
R561 VDPWR.n1550 VDPWR.n163 143.792
R562 VDPWR.n1546 VDPWR.n163 143.792
R563 VDPWR.n981 VDPWR.t31 143.49
R564 VDPWR.n999 VDPWR.t499 143.49
R565 VDPWR.n1017 VDPWR.t6 143.49
R566 VDPWR.n1035 VDPWR.t565 143.49
R567 VDPWR.n1053 VDPWR.t8 143.49
R568 VDPWR.n1071 VDPWR.t142 143.49
R569 VDPWR.n1089 VDPWR.t210 143.49
R570 VDPWR.n1107 VDPWR.t391 143.49
R571 VDPWR.n982 VDPWR.t217 141.511
R572 VDPWR.n1000 VDPWR.t493 141.511
R573 VDPWR.n1018 VDPWR.t279 141.511
R574 VDPWR.n1036 VDPWR.t521 141.511
R575 VDPWR.n1054 VDPWR.t381 141.511
R576 VDPWR.n1072 VDPWR.t104 141.511
R577 VDPWR.n1090 VDPWR.t262 141.511
R578 VDPWR.n1108 VDPWR.t388 141.511
R579 VDPWR.n1538 VDPWR.n1466 139.512
R580 VDPWR.n1512 VDPWR.n1508 139.512
R581 VDPWR.n939 VDPWR.n687 139.512
R582 VDPWR.n846 VDPWR.n841 139.512
R583 VDPWR.n480 VDPWR.n189 139.512
R584 VDPWR.n480 VDPWR.n190 139.512
R585 VDPWR.n484 VDPWR.n183 139.512
R586 VDPWR.n484 VDPWR.n181 139.512
R587 VDPWR.n454 VDPWR.n213 139.512
R588 VDPWR.n454 VDPWR.n214 139.512
R589 VDPWR.n458 VDPWR.n207 139.512
R590 VDPWR.n458 VDPWR.n205 139.512
R591 VDPWR.n428 VDPWR.n237 139.512
R592 VDPWR.n428 VDPWR.n238 139.512
R593 VDPWR.n432 VDPWR.n231 139.512
R594 VDPWR.n432 VDPWR.n229 139.512
R595 VDPWR.n402 VDPWR.n261 139.512
R596 VDPWR.n402 VDPWR.n262 139.512
R597 VDPWR.n406 VDPWR.n255 139.512
R598 VDPWR.n406 VDPWR.n253 139.512
R599 VDPWR.n376 VDPWR.n285 139.512
R600 VDPWR.n376 VDPWR.n286 139.512
R601 VDPWR.n380 VDPWR.n279 139.512
R602 VDPWR.n380 VDPWR.n277 139.512
R603 VDPWR.n342 VDPWR.n309 139.512
R604 VDPWR.n342 VDPWR.n310 139.512
R605 VDPWR.n346 VDPWR.n303 139.512
R606 VDPWR.n346 VDPWR.n301 139.512
R607 VDPWR.n158 VDPWR.n151 139.512
R608 VDPWR.n158 VDPWR.n157 139.512
R609 VDPWR.n111 VDPWR.n20 139.512
R610 VDPWR.n111 VDPWR.n21 139.512
R611 VDPWR.n115 VDPWR.n14 139.512
R612 VDPWR.n115 VDPWR.n12 139.512
R613 VDPWR.n81 VDPWR.n38 139.512
R614 VDPWR.n81 VDPWR.n36 139.512
R615 VDPWR.n77 VDPWR.n45 139.512
R616 VDPWR.n77 VDPWR.n44 139.512
R617 VDPWR.n1172 VDPWR.t227 135.981
R618 VDPWR.n1190 VDPWR.t277 135.981
R619 VDPWR.n1206 VDPWR.t239 135.981
R620 VDPWR.n1222 VDPWR.t85 135.981
R621 VDPWR.n1238 VDPWR.t188 135.981
R622 VDPWR.n1254 VDPWR.t291 135.981
R623 VDPWR.n1270 VDPWR.t57 135.981
R624 VDPWR.n1286 VDPWR.t106 135.981
R625 VDPWR.n1302 VDPWR.t4 135.981
R626 VDPWR.n1373 VDPWR.t16 135.981
R627 VDPWR.t543 VDPWR.n1375 135.981
R628 VDPWR.n1407 VDPWR.t352 135.981
R629 VDPWR.t518 VDPWR.n1401 135.981
R630 VDPWR.n1435 VDPWR.t275 135.981
R631 VDPWR.t126 VDPWR.n1429 135.981
R632 VDPWR.n1459 VDPWR.t299 135.981
R633 VDPWR.n491 VDPWR.n177 135.591
R634 VDPWR.n502 VDPWR.n171 135.591
R635 VDPWR.n130 VDPWR.n8 135.591
R636 VDPWR.n141 VDPWR.n2 135.591
R637 VDPWR.t176 VDPWR.n1173 135.049
R638 VDPWR.t363 VDPWR.n1188 135.049
R639 VDPWR.t256 VDPWR.n1204 135.049
R640 VDPWR.t67 VDPWR.n1220 135.049
R641 VDPWR.t483 VDPWR.n1236 135.049
R642 VDPWR.t393 VDPWR.n1252 135.049
R643 VDPWR.t408 VDPWR.n1268 135.049
R644 VDPWR.t43 VDPWR.n1284 135.049
R645 VDPWR.t224 VDPWR.n1300 135.049
R646 VDPWR.t180 VDPWR.n1378 135.049
R647 VDPWR.n1377 VDPWR.t545 135.049
R648 VDPWR.n1397 VDPWR.t539 135.049
R649 VDPWR.t350 VDPWR.n1399 135.049
R650 VDPWR.t120 VDPWR.n1405 135.049
R651 VDPWR.n1403 VDPWR.t374 135.049
R652 VDPWR.n1425 VDPWR.t379 135.049
R653 VDPWR.t584 VDPWR.n1427 135.049
R654 VDPWR.t212 VDPWR.n1433 135.049
R655 VDPWR.n1431 VDPWR.t87 135.049
R656 VDPWR.n1453 VDPWR.t414 135.049
R657 VDPWR.t53 VDPWR.n1455 135.049
R658 VDPWR.t229 VDPWR.n1457 135.049
R659 VDPWR.n683 VDPWR.n672 134.43
R660 VDPWR.n666 VDPWR.n655 134.43
R661 VDPWR.n649 VDPWR.n638 134.43
R662 VDPWR.n632 VDPWR.n621 134.43
R663 VDPWR.n615 VDPWR.n604 134.43
R664 VDPWR.n598 VDPWR.n587 134.43
R665 VDPWR.n581 VDPWR.n570 134.43
R666 VDPWR.n564 VDPWR.n553 134.43
R667 VDPWR.n1174 VDPWR.t174 132.256
R668 VDPWR.n1189 VDPWR.t570 132.256
R669 VDPWR.n1205 VDPWR.t254 132.256
R670 VDPWR.n1221 VDPWR.t47 132.256
R671 VDPWR.n1237 VDPWR.t476 132.256
R672 VDPWR.n1253 VDPWR.t603 132.256
R673 VDPWR.n1269 VDPWR.t406 132.256
R674 VDPWR.n1285 VDPWR.t45 132.256
R675 VDPWR.n1301 VDPWR.t341 132.256
R676 VDPWR.n1379 VDPWR.t574 132.256
R677 VDPWR.n1374 VDPWR.t233 132.256
R678 VDPWR.n1406 VDPWR.t541 132.256
R679 VDPWR.n1400 VDPWR.t303 132.256
R680 VDPWR.n1434 VDPWR.t39 132.256
R681 VDPWR.n1428 VDPWR.t412 132.256
R682 VDPWR.n1458 VDPWR.t505 132.256
R683 VDPWR.n677 VDPWR.n676 129.874
R684 VDPWR.n676 VDPWR.n672 129.874
R685 VDPWR.n660 VDPWR.n659 129.874
R686 VDPWR.n659 VDPWR.n655 129.874
R687 VDPWR.n643 VDPWR.n642 129.874
R688 VDPWR.n642 VDPWR.n638 129.874
R689 VDPWR.n626 VDPWR.n625 129.874
R690 VDPWR.n625 VDPWR.n621 129.874
R691 VDPWR.n609 VDPWR.n608 129.874
R692 VDPWR.n608 VDPWR.n604 129.874
R693 VDPWR.n592 VDPWR.n591 129.874
R694 VDPWR.n591 VDPWR.n587 129.874
R695 VDPWR.n575 VDPWR.n574 129.874
R696 VDPWR.n574 VDPWR.n570 129.874
R697 VDPWR.n558 VDPWR.n557 129.874
R698 VDPWR.n557 VDPWR.n553 129.874
R699 VDPWR.n496 VDPWR.n175 129.013
R700 VDPWR.n507 VDPWR.n169 129.013
R701 VDPWR.n135 VDPWR.n6 129.013
R702 VDPWR.n146 VDPWR.n0 129.013
R703 VDPWR.n1537 VDPWR.n1469 120.178
R704 VDPWR.n1473 VDPWR.n1471 120.178
R705 VDPWR.n1530 VDPWR.n1476 120.178
R706 VDPWR.n1480 VDPWR.n1478 120.178
R707 VDPWR.n1523 VDPWR.n1483 120.178
R708 VDPWR.n1514 VDPWR.n1513 120.178
R709 VDPWR.n1518 VDPWR.n1485 120.178
R710 VDPWR.n938 VDPWR.n690 120.178
R711 VDPWR.n694 VDPWR.n692 120.178
R712 VDPWR.n931 VDPWR.n697 120.178
R713 VDPWR.n701 VDPWR.n699 120.178
R714 VDPWR.n924 VDPWR.n704 120.178
R715 VDPWR.n708 VDPWR.n706 120.178
R716 VDPWR.n917 VDPWR.n711 120.178
R717 VDPWR.n715 VDPWR.n713 120.178
R718 VDPWR.n910 VDPWR.n718 120.178
R719 VDPWR.n722 VDPWR.n720 120.178
R720 VDPWR.n903 VDPWR.n725 120.178
R721 VDPWR.n729 VDPWR.n727 120.178
R722 VDPWR.n896 VDPWR.n732 120.178
R723 VDPWR.n736 VDPWR.n734 120.178
R724 VDPWR.n889 VDPWR.n739 120.178
R725 VDPWR.n743 VDPWR.n741 120.178
R726 VDPWR.n882 VDPWR.n746 120.178
R727 VDPWR.n750 VDPWR.n748 120.178
R728 VDPWR.n875 VDPWR.n753 120.178
R729 VDPWR.n757 VDPWR.n755 120.178
R730 VDPWR.n868 VDPWR.n760 120.178
R731 VDPWR.n764 VDPWR.n762 120.178
R732 VDPWR.n861 VDPWR.n767 120.178
R733 VDPWR.n771 VDPWR.n769 120.178
R734 VDPWR.n854 VDPWR.n774 120.178
R735 VDPWR.n778 VDPWR.n776 120.178
R736 VDPWR.n847 VDPWR.n781 120.178
R737 VDPWR VDPWR.n1377 108.04
R738 VDPWR.n1399 VDPWR 108.04
R739 VDPWR VDPWR.n1403 108.04
R740 VDPWR.n1427 VDPWR 108.04
R741 VDPWR VDPWR.n1431 108.04
R742 VDPWR.n1455 VDPWR 108.04
R743 VDPWR.t196 VDPWR.t354 88.7478
R744 VDPWR.t418 VDPWR.t199 88.7478
R745 VDPWR.t327 VDPWR.t606 88.7478
R746 VDPWR.t561 VDPWR.t559 88.7478
R747 VDPWR.t163 VDPWR.t165 88.7478
R748 VDPWR.t134 VDPWR.t509 88.7478
R749 VDPWR.t507 VDPWR.t491 88.7478
R750 VDPWR.t130 VDPWR.t426 88.7478
R751 VDPWR.t592 VDPWR.t590 88.7478
R752 VDPWR.t337 VDPWR.t558 88.7478
R753 VDPWR.t243 VDPWR.t171 88.7478
R754 VDPWR.t241 VDPWR.t283 88.7478
R755 VDPWR.t301 VDPWR.t416 88.7478
R756 VDPWR.t285 VDPWR.t226 88.7478
R757 VDPWR.t514 VDPWR.t129 88.7478
R758 VDPWR.t335 VDPWR.t333 88.7478
R759 VDPWR.t610 VDPWR.t97 88.7478
R760 VDPWR.t29 VDPWR.t3 88.7478
R761 VDPWR.t206 VDPWR.t390 88.7478
R762 VDPWR.t220 VDPWR.t208 88.7478
R763 VDPWR.t457 VDPWR.t436 88.7478
R764 VDPWR.t448 VDPWR.t112 88.7478
R765 VDPWR.t512 VDPWR.t520 88.7478
R766 VDPWR.t148 VDPWR.t329 88.7478
R767 VDPWR.t451 VDPWR.t463 88.7478
R768 VDPWR.t439 VDPWR.t511 88.7478
R769 VDPWR.t372 VDPWR.t102 88.7478
R770 VDPWR.t22 VDPWR.t99 88.7478
R771 VDPWR.t460 VDPWR.t433 88.7478
R772 VDPWR.t445 VDPWR.t113 88.7478
R773 VDPWR.t503 VDPWR.t138 88.7478
R774 VDPWR.t501 VDPWR.t582 88.7478
R775 VDPWR.n673 VDPWR.t71 88.2668
R776 VDPWR.n656 VDPWR.t214 88.2668
R777 VDPWR.n639 VDPWR.t315 88.2668
R778 VDPWR.n622 VDPWR.t186 88.2668
R779 VDPWR.n605 VDPWR.t122 88.2668
R780 VDPWR.n588 VDPWR.t246 88.2668
R781 VDPWR.n571 VDPWR.t260 88.2668
R782 VDPWR.n554 VDPWR.t153 88.2668
R783 VDPWR.n675 VDPWR.n673 87.3568
R784 VDPWR.n658 VDPWR.n656 87.3568
R785 VDPWR.n641 VDPWR.n639 87.3568
R786 VDPWR.n624 VDPWR.n622 87.3568
R787 VDPWR.n607 VDPWR.n605 87.3568
R788 VDPWR.n590 VDPWR.n588 87.3568
R789 VDPWR.n573 VDPWR.n571 87.3568
R790 VDPWR.n556 VDPWR.n554 87.3568
R791 VDPWR.t169 VDPWR.t384 87.0838
R792 VDPWR.t33 VDPWR.t169 87.0838
R793 VDPWR.t217 VDPWR.t33 87.0838
R794 VDPWR.t31 VDPWR.t128 87.0838
R795 VDPWR.t128 VDPWR.t497 87.0838
R796 VDPWR.t497 VDPWR.t577 87.0838
R797 VDPWR.t369 VDPWR.t63 87.0838
R798 VDPWR.t533 VDPWR.t369 87.0838
R799 VDPWR.t493 VDPWR.t533 87.0838
R800 VDPWR.t499 VDPWR.t245 87.0838
R801 VDPWR.t245 VDPWR.t580 87.0838
R802 VDPWR.t580 VDPWR.t167 87.0838
R803 VDPWR.t114 VDPWR.t397 87.0838
R804 VDPWR.t266 VDPWR.t114 87.0838
R805 VDPWR.t279 VDPWR.t266 87.0838
R806 VDPWR.t6 VDPWR.t510 87.0838
R807 VDPWR.t510 VDPWR.t399 87.0838
R808 VDPWR.t399 VDPWR.t248 87.0838
R809 VDPWR.t235 VDPWR.t145 87.0838
R810 VDPWR.t264 VDPWR.t235 87.0838
R811 VDPWR.t521 VDPWR.t264 87.0838
R812 VDPWR.t565 VDPWR.t28 87.0838
R813 VDPWR.t28 VDPWR.t356 87.0838
R814 VDPWR.t356 VDPWR.t237 87.0838
R815 VDPWR.t361 VDPWR.t184 87.0838
R816 VDPWR.t84 VDPWR.t361 87.0838
R817 VDPWR.t381 VDPWR.t84 87.0838
R818 VDPWR.t8 VDPWR.t596 87.0838
R819 VDPWR.t596 VDPWR.t182 87.0838
R820 VDPWR.t182 VDPWR.t155 87.0838
R821 VDPWR.t322 VDPWR.t319 87.0838
R822 VDPWR.t125 VDPWR.t322 87.0838
R823 VDPWR.t104 VDPWR.t125 87.0838
R824 VDPWR.t142 VDPWR.t595 87.0838
R825 VDPWR.t595 VDPWR.t317 87.0838
R826 VDPWR.t317 VDPWR.t324 87.0838
R827 VDPWR.t424 VDPWR.t202 87.0838
R828 VDPWR.t101 VDPWR.t424 87.0838
R829 VDPWR.t262 VDPWR.t101 87.0838
R830 VDPWR.t210 VDPWR.t34 87.0838
R831 VDPWR.t34 VDPWR.t204 87.0838
R832 VDPWR.t204 VDPWR.t586 87.0838
R833 VDPWR.t69 VDPWR.t273 87.0838
R834 VDPWR.t468 VDPWR.t69 87.0838
R835 VDPWR.t388 VDPWR.t468 87.0838
R836 VDPWR.t391 VDPWR.t2 87.0838
R837 VDPWR.t2 VDPWR.t345 87.0838
R838 VDPWR.t345 VDPWR.t599 87.0838
R839 VDPWR.n547 VDPWR.t154 85.1439
R840 VDPWR.n542 VDPWR.t532 85.1439
R841 VDPWR.n537 VDPWR.t525 85.1439
R842 VDPWR.n532 VDPWR.t124 85.1439
R843 VDPWR.n527 VDPWR.t259 85.1439
R844 VDPWR.n522 VDPWR.t488 85.1439
R845 VDPWR.n517 VDPWR.t258 85.1439
R846 VDPWR.n512 VDPWR.t401 85.1439
R847 VDPWR.n973 VDPWR.t218 85.0216
R848 VDPWR.n988 VDPWR.t32 85.0216
R849 VDPWR.n969 VDPWR.t494 85.0216
R850 VDPWR.n1006 VDPWR.t500 85.0216
R851 VDPWR.n965 VDPWR.t280 85.0216
R852 VDPWR.n1024 VDPWR.t7 85.0216
R853 VDPWR.n961 VDPWR.t522 85.0216
R854 VDPWR.n1042 VDPWR.t566 85.0216
R855 VDPWR.n957 VDPWR.t382 85.0216
R856 VDPWR.n1060 VDPWR.t9 85.0216
R857 VDPWR.n953 VDPWR.t105 85.0216
R858 VDPWR.n1078 VDPWR.t143 85.0216
R859 VDPWR.n949 VDPWR.t263 85.0216
R860 VDPWR.n1096 VDPWR.t211 85.0216
R861 VDPWR.n945 VDPWR.t389 85.0216
R862 VDPWR.n1114 VDPWR.t392 85.0216
R863 VDPWR.n166 VDPWR.t140 84.9265
R864 VDPWR.n162 VDPWR.t534 84.9265
R865 VDPWR.n1510 VDPWR.t469 84.9238
R866 VDPWR.n1503 VDPWR.t161 84.9238
R867 VDPWR.n48 VDPWR.n47 84.8474
R868 VDPWR.n1467 VDPWR.t83 84.7934
R869 VDPWR.n1534 VDPWR.t198 84.7934
R870 VDPWR.n1474 VDPWR.t326 84.7934
R871 VDPWR.n1527 VDPWR.t160 84.7934
R872 VDPWR.n1481 VDPWR.t162 84.7934
R873 VDPWR.n1520 VDPWR.t159 84.7934
R874 VDPWR.n688 VDPWR.t607 84.7934
R875 VDPWR.n935 VDPWR.t150 84.7934
R876 VDPWR.n695 VDPWR.t110 84.7934
R877 VDPWR.n928 VDPWR.t147 84.7934
R878 VDPWR.n702 VDPWR.t405 84.7934
R879 VDPWR.n921 VDPWR.t193 84.7934
R880 VDPWR.n709 VDPWR.t609 84.7934
R881 VDPWR.n914 VDPWR.t404 84.7934
R882 VDPWR.n716 VDPWR.t173 84.7934
R883 VDPWR.n907 VDPWR.t602 84.7934
R884 VDPWR.n723 VDPWR.t172 84.7934
R885 VDPWR.n900 VDPWR.t601 84.7934
R886 VDPWR.n730 VDPWR.t192 84.7934
R887 VDPWR.n893 VDPWR.t608 84.7934
R888 VDPWR.n737 VDPWR.t403 84.7934
R889 VDPWR.n886 VDPWR.t111 84.7934
R890 VDPWR.n744 VDPWR.t554 84.7934
R891 VDPWR.n879 VDPWR.t556 84.7934
R892 VDPWR.n751 VDPWR.t557 84.7934
R893 VDPWR.n872 VDPWR.t555 84.7934
R894 VDPWR.n758 VDPWR.t25 84.7934
R895 VDPWR.n865 VDPWR.t482 84.7934
R896 VDPWR.n765 VDPWR.t103 84.7934
R897 VDPWR.n858 VDPWR.t594 84.7934
R898 VDPWR.n772 VDPWR.t265 84.7934
R899 VDPWR.n851 VDPWR.t597 84.7934
R900 VDPWR.n779 VDPWR.t81 84.7934
R901 VDPWR.n844 VDPWR.t141 84.7934
R902 VDPWR.n478 VDPWR.t589 84.7934
R903 VDPWR.n486 VDPWR.t340 84.7934
R904 VDPWR.n452 VDPWR.t605 84.7934
R905 VDPWR.n460 VDPWR.t137 84.7934
R906 VDPWR.n426 VDPWR.t387 84.7934
R907 VDPWR.n434 VDPWR.t567 84.7934
R908 VDPWR.n400 VDPWR.t251 84.7934
R909 VDPWR.n408 VDPWR.t553 84.7934
R910 VDPWR.n374 VDPWR.t368 84.7934
R911 VDPWR.n382 VDPWR.t612 84.7934
R912 VDPWR.n340 VDPWR.t579 84.7934
R913 VDPWR.n348 VDPWR.t467 84.7934
R914 VDPWR.n152 VDPWR.t332 84.7934
R915 VDPWR.n109 VDPWR.t485 84.7934
R916 VDPWR.n117 VDPWR.t443 84.7934
R917 VDPWR.n75 VDPWR.t598 84.7934
R918 VDPWR.n83 VDPWR.t455 84.7934
R919 VDPWR.n549 VDPWR.t588 84.7906
R920 VDPWR.n547 VDPWR.t383 84.7906
R921 VDPWR.n548 VDPWR.t576 84.7906
R922 VDPWR.n544 VDPWR.t402 84.7906
R923 VDPWR.n542 VDPWR.t261 84.7906
R924 VDPWR.n543 VDPWR.t371 84.7906
R925 VDPWR.n539 VDPWR.t492 84.7906
R926 VDPWR.n537 VDPWR.t479 84.7906
R927 VDPWR.n538 VDPWR.t247 84.7906
R928 VDPWR.n534 VDPWR.t216 84.7906
R929 VDPWR.n532 VDPWR.t144 84.7906
R930 VDPWR.n533 VDPWR.t123 84.7906
R931 VDPWR.n529 VDPWR.t489 84.7906
R932 VDPWR.n527 VDPWR.t187 84.7906
R933 VDPWR.n528 VDPWR.t360 84.7906
R934 VDPWR.n524 VDPWR.t378 84.7906
R935 VDPWR.n522 VDPWR.t316 84.7906
R936 VDPWR.n523 VDPWR.t321 84.7906
R937 VDPWR.n519 VDPWR.t215 84.7906
R938 VDPWR.n517 VDPWR.t219 84.7906
R939 VDPWR.n518 VDPWR.t478 84.7906
R940 VDPWR.n514 VDPWR.t490 84.7906
R941 VDPWR.n512 VDPWR.t347 84.7906
R942 VDPWR.n513 VDPWR.t72 84.7906
R943 VDPWR.n489 VDPWR.t223 84.7771
R944 VDPWR.n500 VDPWR.t179 84.7771
R945 VDPWR.n128 VDPWR.t78 84.7771
R946 VDPWR.n139 VDPWR.t473 84.7771
R947 VDPWR.n204 VDPWR.n203 84.7744
R948 VDPWR.n193 VDPWR.n192 84.7744
R949 VDPWR.n228 VDPWR.n227 84.7744
R950 VDPWR.n217 VDPWR.n216 84.7744
R951 VDPWR.n252 VDPWR.n251 84.7744
R952 VDPWR.n241 VDPWR.n240 84.7744
R953 VDPWR.n276 VDPWR.n275 84.7744
R954 VDPWR.n265 VDPWR.n264 84.7744
R955 VDPWR.n300 VDPWR.n299 84.7744
R956 VDPWR.n289 VDPWR.n288 84.7744
R957 VDPWR.n324 VDPWR.n323 84.7744
R958 VDPWR.n313 VDPWR.n312 84.7744
R959 VDPWR.n35 VDPWR.n34 84.7744
R960 VDPWR.n24 VDPWR.n23 84.7744
R961 VDPWR.n59 VDPWR.n58 84.7744
R962 VDPWR.n498 VDPWR.t21 84.7716
R963 VDPWR.n509 VDPWR.t1 84.7716
R964 VDPWR.n137 VDPWR.t573 84.7716
R965 VDPWR.n148 VDPWR.t27 84.7716
R966 VDPWR.n204 VDPWR.t197 83.8097
R967 VDPWR.n193 VDPWR.t560 83.8097
R968 VDPWR.n228 VDPWR.t164 83.8097
R969 VDPWR.n217 VDPWR.t427 83.8097
R970 VDPWR.n252 VDPWR.t593 83.8097
R971 VDPWR.n241 VDPWR.t284 83.8097
R972 VDPWR.n276 VDPWR.t302 83.8097
R973 VDPWR.n265 VDPWR.t334 83.8097
R974 VDPWR.n300 VDPWR.t611 83.8097
R975 VDPWR.n289 VDPWR.t209 83.8097
R976 VDPWR.n324 VDPWR.t458 83.8097
R977 VDPWR.n313 VDPWR.t330 83.8097
R978 VDPWR.n35 VDPWR.t452 83.8097
R979 VDPWR.n24 VDPWR.t100 83.8097
R980 VDPWR.n59 VDPWR.t461 83.8097
R981 VDPWR.n48 VDPWR.t583 83.8097
R982 VDPWR.t535 VDPWR.t470 81.9613
R983 VDPWR.t132 VDPWR.t535 81.9613
R984 VDPWR.t227 VDPWR.t132 81.9613
R985 VDPWR.t174 VDPWR.t35 81.9613
R986 VDPWR.t35 VDPWR.t348 81.9613
R987 VDPWR.t348 VDPWR.t176 81.9613
R988 VDPWR.t551 VDPWR.t547 81.9613
R989 VDPWR.t549 VDPWR.t551 81.9613
R990 VDPWR.t277 VDPWR.t549 81.9613
R991 VDPWR.t570 VDPWR.t568 81.9613
R992 VDPWR.t568 VDPWR.t523 81.9613
R993 VDPWR.t523 VDPWR.t363 81.9613
R994 VDPWR.t516 VDPWR.t194 81.9613
R995 VDPWR.t376 VDPWR.t516 81.9613
R996 VDPWR.t239 VDPWR.t376 81.9613
R997 VDPWR.t254 VDPWR.t311 81.9613
R998 VDPWR.t311 VDPWR.t309 81.9613
R999 VDPWR.t309 VDPWR.t256 81.9613
R1000 VDPWR.t537 VDPWR.t61 81.9613
R1001 VDPWR.t231 VDPWR.t537 81.9613
R1002 VDPWR.t85 VDPWR.t231 81.9613
R1003 VDPWR.t47 VDPWR.t495 81.9613
R1004 VDPWR.t495 VDPWR.t79 81.9613
R1005 VDPWR.t79 VDPWR.t67 81.9613
R1006 VDPWR.t41 VDPWR.t281 81.9613
R1007 VDPWR.t190 VDPWR.t41 81.9613
R1008 VDPWR.t188 VDPWR.t190 81.9613
R1009 VDPWR.t476 VDPWR.t474 81.9613
R1010 VDPWR.t474 VDPWR.t297 81.9613
R1011 VDPWR.t297 VDPWR.t483 81.9613
R1012 VDPWR.t287 VDPWR.t293 81.9613
R1013 VDPWR.t289 VDPWR.t287 81.9613
R1014 VDPWR.t291 VDPWR.t289 81.9613
R1015 VDPWR.t603 VDPWR.t395 81.9613
R1016 VDPWR.t395 VDPWR.t295 81.9613
R1017 VDPWR.t295 VDPWR.t393 81.9613
R1018 VDPWR.t118 VDPWR.t526 81.9613
R1019 VDPWR.t59 VDPWR.t118 81.9613
R1020 VDPWR.t57 VDPWR.t59 81.9613
R1021 VDPWR.t406 VDPWR.t410 81.9613
R1022 VDPWR.t410 VDPWR.t430 81.9613
R1023 VDPWR.t430 VDPWR.t408 81.9613
R1024 VDPWR.t37 VDPWR.t108 81.9613
R1025 VDPWR.t428 VDPWR.t37 81.9613
R1026 VDPWR.t106 VDPWR.t428 81.9613
R1027 VDPWR.t45 VDPWR.t528 81.9613
R1028 VDPWR.t528 VDPWR.t613 81.9613
R1029 VDPWR.t613 VDPWR.t43 81.9613
R1030 VDPWR.t563 VDPWR.t12 81.9613
R1031 VDPWR.t10 VDPWR.t563 81.9613
R1032 VDPWR.t4 VDPWR.t10 81.9613
R1033 VDPWR.t341 VDPWR.t267 81.9613
R1034 VDPWR.t267 VDPWR.t65 81.9613
R1035 VDPWR.t65 VDPWR.t224 81.9613
R1036 VDPWR.t93 VDPWR.t14 81.9613
R1037 VDPWR.t18 VDPWR.t93 81.9613
R1038 VDPWR.t16 VDPWR.t18 81.9613
R1039 VDPWR.t574 VDPWR.t51 81.9613
R1040 VDPWR.t51 VDPWR.t358 81.9613
R1041 VDPWR.t358 VDPWR.t180 81.9613
R1042 VDPWR.t545 VDPWR.t269 81.9613
R1043 VDPWR.t269 VDPWR.t252 81.9613
R1044 VDPWR.t252 VDPWR.t543 81.9613
R1045 VDPWR.t233 VDPWR.t55 81.9613
R1046 VDPWR.t55 VDPWR.t116 81.9613
R1047 VDPWR.t116 VDPWR.t539 81.9613
R1048 VDPWR.t486 VDPWR.t350 81.9613
R1049 VDPWR.t480 VDPWR.t486 81.9613
R1050 VDPWR.t352 VDPWR.t480 81.9613
R1051 VDPWR.t541 VDPWR.t157 81.9613
R1052 VDPWR.t157 VDPWR.t151 81.9613
R1053 VDPWR.t151 VDPWR.t120 81.9613
R1054 VDPWR.t374 VDPWR.t530 81.9613
R1055 VDPWR.t530 VDPWR.t75 81.9613
R1056 VDPWR.t75 VDPWR.t518 81.9613
R1057 VDPWR.t303 VDPWR.t307 81.9613
R1058 VDPWR.t307 VDPWR.t305 81.9613
R1059 VDPWR.t305 VDPWR.t379 81.9613
R1060 VDPWR.t271 VDPWR.t584 81.9613
R1061 VDPWR.t343 VDPWR.t271 81.9613
R1062 VDPWR.t275 VDPWR.t343 81.9613
R1063 VDPWR.t39 VDPWR.t95 81.9613
R1064 VDPWR.t95 VDPWR.t313 81.9613
R1065 VDPWR.t313 VDPWR.t212 81.9613
R1066 VDPWR.t87 VDPWR.t365 81.9613
R1067 VDPWR.t365 VDPWR.t73 81.9613
R1068 VDPWR.t73 VDPWR.t126 81.9613
R1069 VDPWR.t412 VDPWR.t91 81.9613
R1070 VDPWR.t91 VDPWR.t89 81.9613
R1071 VDPWR.t89 VDPWR.t414 81.9613
R1072 VDPWR.t422 VDPWR.t53 81.9613
R1073 VDPWR.t420 VDPWR.t422 81.9613
R1074 VDPWR.t299 VDPWR.t420 81.9613
R1075 VDPWR.t505 VDPWR.t49 81.9613
R1076 VDPWR.t49 VDPWR.t200 81.9613
R1077 VDPWR.t200 VDPWR.t229 81.9613
R1078 VDPWR.n1368 VDPWR.n1367 75.8478
R1079 VDPWR.n1363 VDPWR.n1362 75.7173
R1080 VDPWR.n1383 VDPWR.n1361 75.7173
R1081 VDPWR.n1384 VDPWR.n1360 75.7173
R1082 VDPWR.n1387 VDPWR.n1358 75.7173
R1083 VDPWR.n1388 VDPWR.n1357 75.7173
R1084 VDPWR.n1392 VDPWR.n1389 75.7173
R1085 VDPWR.n1391 VDPWR.n1390 75.7173
R1086 VDPWR.n1352 VDPWR.n1351 75.7173
R1087 VDPWR.n1347 VDPWR.n1346 75.7173
R1088 VDPWR.n1411 VDPWR.n1345 75.7173
R1089 VDPWR.n1412 VDPWR.n1344 75.7173
R1090 VDPWR.n1415 VDPWR.n1342 75.7173
R1091 VDPWR.n1416 VDPWR.n1341 75.7173
R1092 VDPWR.n1420 VDPWR.n1417 75.7173
R1093 VDPWR.n1419 VDPWR.n1418 75.7173
R1094 VDPWR.n1336 VDPWR.n1335 75.7173
R1095 VDPWR.n1331 VDPWR.n1330 75.7173
R1096 VDPWR.n1439 VDPWR.n1329 75.7173
R1097 VDPWR.n1440 VDPWR.n1328 75.7173
R1098 VDPWR.n1443 VDPWR.n1326 75.7173
R1099 VDPWR.n1444 VDPWR.n1325 75.7173
R1100 VDPWR.n1448 VDPWR.n1445 75.7173
R1101 VDPWR.n1447 VDPWR.n1446 75.7173
R1102 VDPWR.n1320 VDPWR.n1319 75.7173
R1103 VDPWR.n1315 VDPWR.n1314 75.7173
R1104 VDPWR.n1463 VDPWR.n1313 75.7173
R1105 VDPWR.n1464 VDPWR.n1312 75.7173
R1106 VDPWR.n1168 VDPWR.n1167 75.7173
R1107 VDPWR.n1163 VDPWR.n1162 75.7173
R1108 VDPWR.n1178 VDPWR.n1161 75.7173
R1109 VDPWR.n1179 VDPWR.n1160 75.7173
R1110 VDPWR.n1182 VDPWR.n1181 75.7173
R1111 VDPWR.n1158 VDPWR.n1157 75.7173
R1112 VDPWR.n1194 VDPWR.n1156 75.7173
R1113 VDPWR.n1195 VDPWR.n1155 75.7173
R1114 VDPWR.n1198 VDPWR.n1197 75.7173
R1115 VDPWR.n1153 VDPWR.n1152 75.7173
R1116 VDPWR.n1210 VDPWR.n1151 75.7173
R1117 VDPWR.n1211 VDPWR.n1150 75.7173
R1118 VDPWR.n1214 VDPWR.n1213 75.7173
R1119 VDPWR.n1148 VDPWR.n1147 75.7173
R1120 VDPWR.n1226 VDPWR.n1146 75.7173
R1121 VDPWR.n1227 VDPWR.n1145 75.7173
R1122 VDPWR.n1230 VDPWR.n1229 75.7173
R1123 VDPWR.n1143 VDPWR.n1142 75.7173
R1124 VDPWR.n1242 VDPWR.n1141 75.7173
R1125 VDPWR.n1243 VDPWR.n1140 75.7173
R1126 VDPWR.n1246 VDPWR.n1245 75.7173
R1127 VDPWR.n1138 VDPWR.n1137 75.7173
R1128 VDPWR.n1258 VDPWR.n1136 75.7173
R1129 VDPWR.n1259 VDPWR.n1135 75.7173
R1130 VDPWR.n1262 VDPWR.n1261 75.7173
R1131 VDPWR.n1133 VDPWR.n1132 75.7173
R1132 VDPWR.n1274 VDPWR.n1131 75.7173
R1133 VDPWR.n1275 VDPWR.n1130 75.7173
R1134 VDPWR.n1278 VDPWR.n1277 75.7173
R1135 VDPWR.n1128 VDPWR.n1127 75.7173
R1136 VDPWR.n1290 VDPWR.n1126 75.7173
R1137 VDPWR.n1291 VDPWR.n1125 75.7173
R1138 VDPWR.n1294 VDPWR.n1293 75.7173
R1139 VDPWR.n1123 VDPWR.n1122 75.7173
R1140 VDPWR.n1306 VDPWR.n1121 75.7173
R1141 VDPWR.n1307 VDPWR.n1120 75.7173
R1142 VDPWR.n975 VDPWR.n974 75.5
R1143 VDPWR.n989 VDPWR.n971 75.5
R1144 VDPWR.n992 VDPWR.n991 75.5
R1145 VDPWR.n1007 VDPWR.n967 75.5
R1146 VDPWR.n1010 VDPWR.n1009 75.5
R1147 VDPWR.n1025 VDPWR.n963 75.5
R1148 VDPWR.n1028 VDPWR.n1027 75.5
R1149 VDPWR.n1043 VDPWR.n959 75.5
R1150 VDPWR.n1046 VDPWR.n1045 75.5
R1151 VDPWR.n1061 VDPWR.n955 75.5
R1152 VDPWR.n1064 VDPWR.n1063 75.5
R1153 VDPWR.n1079 VDPWR.n951 75.5
R1154 VDPWR.n1082 VDPWR.n1081 75.5
R1155 VDPWR.n1097 VDPWR.n947 75.5
R1156 VDPWR.n1100 VDPWR.n1099 75.5
R1157 VDPWR.n1115 VDPWR.n943 75.5
R1158 VDPWR.n495 VDPWR.n178 61.6672
R1159 VDPWR.n506 VDPWR.n172 61.6672
R1160 VDPWR.n134 VDPWR.n9 61.6672
R1161 VDPWR.n145 VDPWR.n3 61.6672
R1162 VDPWR.n155 VDPWR.t331 57.2869
R1163 VDPWR.n1173 VDPWR 50.2946
R1164 VDPWR.n1188 VDPWR 50.2946
R1165 VDPWR.n1204 VDPWR 50.2946
R1166 VDPWR.n1220 VDPWR 50.2946
R1167 VDPWR.n1236 VDPWR 50.2946
R1168 VDPWR.n1252 VDPWR 50.2946
R1169 VDPWR.n1268 VDPWR 50.2946
R1170 VDPWR.n1284 VDPWR 50.2946
R1171 VDPWR.n1300 VDPWR 50.2946
R1172 VDPWR.n1378 VDPWR 50.2946
R1173 VDPWR VDPWR.n1397 50.2946
R1174 VDPWR.n1405 VDPWR 50.2946
R1175 VDPWR VDPWR.n1425 50.2946
R1176 VDPWR.n1433 VDPWR 50.2946
R1177 VDPWR VDPWR.n1453 50.2946
R1178 VDPWR.n1457 VDPWR 50.2946
R1179 VDPWR.n1512 VDPWR.n1507 46.2505
R1180 VDPWR.n1507 VDPWR.n1501 46.2505
R1181 VDPWR.n1506 VDPWR.n1505 46.2505
R1182 VDPWR.n1505 VDPWR.n1501 46.2505
R1183 VDPWR.n1522 VDPWR.n1484 46.2505
R1184 VDPWR.n1501 VDPWR.n1484 46.2505
R1185 VDPWR.n1524 VDPWR.n1482 46.2505
R1186 VDPWR.n1501 VDPWR.n1482 46.2505
R1187 VDPWR.n1529 VDPWR.n1477 46.2505
R1188 VDPWR.n1501 VDPWR.n1477 46.2505
R1189 VDPWR.n1531 VDPWR.n1475 46.2505
R1190 VDPWR.n1501 VDPWR.n1475 46.2505
R1191 VDPWR.n1536 VDPWR.n1470 46.2505
R1192 VDPWR.n1501 VDPWR.n1470 46.2505
R1193 VDPWR.n1538 VDPWR.n1468 46.2505
R1194 VDPWR.n1501 VDPWR.n1468 46.2505
R1195 VDPWR.n846 VDPWR.n782 46.2505
R1196 VDPWR.n836 VDPWR.n782 46.2505
R1197 VDPWR.n848 VDPWR.n780 46.2505
R1198 VDPWR.n836 VDPWR.n780 46.2505
R1199 VDPWR.n853 VDPWR.n775 46.2505
R1200 VDPWR.n836 VDPWR.n775 46.2505
R1201 VDPWR.n855 VDPWR.n773 46.2505
R1202 VDPWR.n836 VDPWR.n773 46.2505
R1203 VDPWR.n860 VDPWR.n768 46.2505
R1204 VDPWR.n836 VDPWR.n768 46.2505
R1205 VDPWR.n862 VDPWR.n766 46.2505
R1206 VDPWR.n836 VDPWR.n766 46.2505
R1207 VDPWR.n867 VDPWR.n761 46.2505
R1208 VDPWR.n836 VDPWR.n761 46.2505
R1209 VDPWR.n869 VDPWR.n759 46.2505
R1210 VDPWR.n836 VDPWR.n759 46.2505
R1211 VDPWR.n874 VDPWR.n754 46.2505
R1212 VDPWR.n836 VDPWR.n754 46.2505
R1213 VDPWR.n876 VDPWR.n752 46.2505
R1214 VDPWR.n836 VDPWR.n752 46.2505
R1215 VDPWR.n881 VDPWR.n747 46.2505
R1216 VDPWR.n836 VDPWR.n747 46.2505
R1217 VDPWR.n883 VDPWR.n745 46.2505
R1218 VDPWR.n836 VDPWR.n745 46.2505
R1219 VDPWR.n888 VDPWR.n740 46.2505
R1220 VDPWR.n836 VDPWR.n740 46.2505
R1221 VDPWR.n890 VDPWR.n738 46.2505
R1222 VDPWR.n836 VDPWR.n738 46.2505
R1223 VDPWR.n895 VDPWR.n733 46.2505
R1224 VDPWR.n836 VDPWR.n733 46.2505
R1225 VDPWR.n897 VDPWR.n731 46.2505
R1226 VDPWR.n836 VDPWR.n731 46.2505
R1227 VDPWR.n902 VDPWR.n726 46.2505
R1228 VDPWR.n836 VDPWR.n726 46.2505
R1229 VDPWR.n904 VDPWR.n724 46.2505
R1230 VDPWR.n836 VDPWR.n724 46.2505
R1231 VDPWR.n909 VDPWR.n719 46.2505
R1232 VDPWR.n836 VDPWR.n719 46.2505
R1233 VDPWR.n911 VDPWR.n717 46.2505
R1234 VDPWR.n836 VDPWR.n717 46.2505
R1235 VDPWR.n916 VDPWR.n712 46.2505
R1236 VDPWR.n836 VDPWR.n712 46.2505
R1237 VDPWR.n918 VDPWR.n710 46.2505
R1238 VDPWR.n836 VDPWR.n710 46.2505
R1239 VDPWR.n923 VDPWR.n705 46.2505
R1240 VDPWR.n836 VDPWR.n705 46.2505
R1241 VDPWR.n925 VDPWR.n703 46.2505
R1242 VDPWR.n836 VDPWR.n703 46.2505
R1243 VDPWR.n930 VDPWR.n698 46.2505
R1244 VDPWR.n836 VDPWR.n698 46.2505
R1245 VDPWR.n932 VDPWR.n696 46.2505
R1246 VDPWR.n836 VDPWR.n696 46.2505
R1247 VDPWR.n937 VDPWR.n691 46.2505
R1248 VDPWR.n836 VDPWR.n691 46.2505
R1249 VDPWR.n939 VDPWR.n689 46.2505
R1250 VDPWR.n836 VDPWR.n689 46.2505
R1251 VDPWR.n481 VDPWR.n480 46.2505
R1252 VDPWR.n482 VDPWR.n481 46.2505
R1253 VDPWR.n484 VDPWR.n483 46.2505
R1254 VDPWR.n483 VDPWR.n482 46.2505
R1255 VDPWR.n455 VDPWR.n454 46.2505
R1256 VDPWR.n456 VDPWR.n455 46.2505
R1257 VDPWR.n458 VDPWR.n457 46.2505
R1258 VDPWR.n457 VDPWR.n456 46.2505
R1259 VDPWR.n429 VDPWR.n428 46.2505
R1260 VDPWR.n430 VDPWR.n429 46.2505
R1261 VDPWR.n432 VDPWR.n431 46.2505
R1262 VDPWR.n431 VDPWR.n430 46.2505
R1263 VDPWR.n403 VDPWR.n402 46.2505
R1264 VDPWR.n404 VDPWR.n403 46.2505
R1265 VDPWR.n406 VDPWR.n405 46.2505
R1266 VDPWR.n405 VDPWR.n404 46.2505
R1267 VDPWR.n377 VDPWR.n376 46.2505
R1268 VDPWR.n378 VDPWR.n377 46.2505
R1269 VDPWR.n380 VDPWR.n379 46.2505
R1270 VDPWR.n379 VDPWR.n378 46.2505
R1271 VDPWR.n343 VDPWR.n342 46.2505
R1272 VDPWR.n344 VDPWR.n343 46.2505
R1273 VDPWR.n346 VDPWR.n345 46.2505
R1274 VDPWR.n345 VDPWR.n344 46.2505
R1275 VDPWR.n158 VDPWR.n153 46.2505
R1276 VDPWR.n112 VDPWR.n111 46.2505
R1277 VDPWR.n113 VDPWR.n112 46.2505
R1278 VDPWR.n115 VDPWR.n114 46.2505
R1279 VDPWR.n114 VDPWR.n113 46.2505
R1280 VDPWR.n81 VDPWR.n80 46.2505
R1281 VDPWR.n80 VDPWR.n79 46.2505
R1282 VDPWR.n78 VDPWR.n77 46.2505
R1283 VDPWR.n79 VDPWR.n78 46.2505
R1284 VDPWR.n1548 VDPWR.t139 44.5923
R1285 VDPWR.n839 VDPWR.n836 44.5678
R1286 VDPWR.t354 VDPWR.n200 44.3742
R1287 VDPWR.n200 VDPWR.t418 44.3742
R1288 VDPWR.n470 VDPWR.t327 44.3742
R1289 VDPWR.n470 VDPWR.t561 44.3742
R1290 VDPWR.t165 VDPWR.n224 44.3742
R1291 VDPWR.n224 VDPWR.t134 44.3742
R1292 VDPWR.n444 VDPWR.t507 44.3742
R1293 VDPWR.n444 VDPWR.t130 44.3742
R1294 VDPWR.t590 VDPWR.n248 44.3742
R1295 VDPWR.n248 VDPWR.t337 44.3742
R1296 VDPWR.n418 VDPWR.t243 44.3742
R1297 VDPWR.n418 VDPWR.t241 44.3742
R1298 VDPWR.t416 VDPWR.n272 44.3742
R1299 VDPWR.n272 VDPWR.t285 44.3742
R1300 VDPWR.n392 VDPWR.t514 44.3742
R1301 VDPWR.n392 VDPWR.t335 44.3742
R1302 VDPWR.t97 VDPWR.n296 44.3742
R1303 VDPWR.n296 VDPWR.t29 44.3742
R1304 VDPWR.n366 VDPWR.t206 44.3742
R1305 VDPWR.n366 VDPWR.t220 44.3742
R1306 VDPWR.t436 VDPWR.n320 44.3742
R1307 VDPWR.n320 VDPWR.t448 44.3742
R1308 VDPWR.n332 VDPWR.t512 44.3742
R1309 VDPWR.n332 VDPWR.t148 44.3742
R1310 VDPWR.t463 VDPWR.n31 44.3742
R1311 VDPWR.n31 VDPWR.t439 44.3742
R1312 VDPWR.n101 VDPWR.t372 44.3742
R1313 VDPWR.n101 VDPWR.t22 44.3742
R1314 VDPWR.t433 VDPWR.n55 44.3742
R1315 VDPWR.n55 VDPWR.t445 44.3742
R1316 VDPWR.n67 VDPWR.t503 44.3742
R1317 VDPWR.n67 VDPWR.t501 44.3742
R1318 VDPWR.n179 VDPWR.n177 43.625
R1319 VDPWR.n173 VDPWR.n171 43.625
R1320 VDPWR.n10 VDPWR.n8 43.625
R1321 VDPWR.n4 VDPWR.n2 43.625
R1322 VDPWR.n505 VDPWR.n169 35.5442
R1323 VDPWR.n144 VDPWR.n0 35.5442
R1324 VDPWR.n494 VDPWR.n175 35.5275
R1325 VDPWR.n133 VDPWR.n6 35.5275
R1326 VDPWR.n1547 VDPWR.n1546 33.509
R1327 VDPWR.n157 VDPWR.n156 32.2656
R1328 VDPWR.n555 VDPWR.n552 31.5192
R1329 VDPWR.n572 VDPWR.n569 31.5192
R1330 VDPWR.n589 VDPWR.n586 31.5192
R1331 VDPWR.n606 VDPWR.n603 31.5192
R1332 VDPWR.n623 VDPWR.n620 31.5192
R1333 VDPWR.n640 VDPWR.n637 31.5192
R1334 VDPWR.n657 VDPWR.n654 31.5192
R1335 VDPWR.n674 VDPWR.n671 31.5192
R1336 VDPWR.n186 VDPWR.t339 28.6437
R1337 VDPWR.n210 VDPWR.t136 28.6437
R1338 VDPWR.n234 VDPWR.t386 28.6437
R1339 VDPWR.n258 VDPWR.t250 28.6437
R1340 VDPWR.n282 VDPWR.t367 28.6437
R1341 VDPWR.n306 VDPWR.t466 28.6437
R1342 VDPWR.n17 VDPWR.t442 28.6437
R1343 VDPWR.n41 VDPWR.t454 28.6437
R1344 VDPWR.n465 VDPWR.n198 23.1255
R1345 VDPWR.n200 VDPWR.n198 23.1255
R1346 VDPWR.n472 VDPWR.n471 23.1255
R1347 VDPWR.n471 VDPWR.n470 23.1255
R1348 VDPWR.n439 VDPWR.n222 23.1255
R1349 VDPWR.n224 VDPWR.n222 23.1255
R1350 VDPWR.n446 VDPWR.n445 23.1255
R1351 VDPWR.n445 VDPWR.n444 23.1255
R1352 VDPWR.n413 VDPWR.n246 23.1255
R1353 VDPWR.n248 VDPWR.n246 23.1255
R1354 VDPWR.n420 VDPWR.n419 23.1255
R1355 VDPWR.n419 VDPWR.n418 23.1255
R1356 VDPWR.n387 VDPWR.n270 23.1255
R1357 VDPWR.n272 VDPWR.n270 23.1255
R1358 VDPWR.n394 VDPWR.n393 23.1255
R1359 VDPWR.n393 VDPWR.n392 23.1255
R1360 VDPWR.n361 VDPWR.n294 23.1255
R1361 VDPWR.n296 VDPWR.n294 23.1255
R1362 VDPWR.n368 VDPWR.n367 23.1255
R1363 VDPWR.n367 VDPWR.n366 23.1255
R1364 VDPWR.n327 VDPWR.n318 23.1255
R1365 VDPWR.n320 VDPWR.n318 23.1255
R1366 VDPWR.n334 VDPWR.n333 23.1255
R1367 VDPWR.n333 VDPWR.n332 23.1255
R1368 VDPWR.n96 VDPWR.n29 23.1255
R1369 VDPWR.n31 VDPWR.n29 23.1255
R1370 VDPWR.n103 VDPWR.n102 23.1255
R1371 VDPWR.n102 VDPWR.n101 23.1255
R1372 VDPWR.n62 VDPWR.n53 23.1255
R1373 VDPWR.n55 VDPWR.n53 23.1255
R1374 VDPWR.n69 VDPWR.n68 23.1255
R1375 VDPWR.n68 VDPWR.n67 23.1255
R1376 VDPWR.n493 VDPWR.t20 20.8338
R1377 VDPWR.n132 VDPWR.t572 20.8338
R1378 VDPWR.n504 VDPWR.t0 20.7429
R1379 VDPWR.n143 VDPWR.t26 20.7429
R1380 VDPWR.n1499 VDPWR.n1483 20.5561
R1381 VDPWR.n1516 VDPWR.n1499 20.5561
R1382 VDPWR.n1497 VDPWR.n1480 20.5561
R1383 VDPWR.n1516 VDPWR.n1497 20.5561
R1384 VDPWR.n1495 VDPWR.n1476 20.5561
R1385 VDPWR.n1516 VDPWR.n1495 20.5561
R1386 VDPWR.n1493 VDPWR.n1473 20.5561
R1387 VDPWR.n1516 VDPWR.n1493 20.5561
R1388 VDPWR.n1491 VDPWR.n1469 20.5561
R1389 VDPWR.n1516 VDPWR.n1491 20.5561
R1390 VDPWR.n1489 VDPWR.n1466 20.5561
R1391 VDPWR.n1516 VDPWR.n1489 20.5561
R1392 VDPWR.n1515 VDPWR.n1514 20.5561
R1393 VDPWR.n1516 VDPWR.n1515 20.5561
R1394 VDPWR.n1508 VDPWR.n1500 20.5561
R1395 VDPWR.n1516 VDPWR.n1500 20.5561
R1396 VDPWR.n1518 VDPWR.n1517 20.5561
R1397 VDPWR.n1517 VDPWR.n1516 20.5561
R1398 VDPWR.n977 VDPWR.n976 20.5561
R1399 VDPWR.n980 VDPWR.n972 20.5561
R1400 VDPWR.n981 VDPWR.n980 20.5561
R1401 VDPWR.n979 VDPWR.n970 20.5561
R1402 VDPWR.n995 VDPWR.n994 20.5561
R1403 VDPWR.n998 VDPWR.n968 20.5561
R1404 VDPWR.n999 VDPWR.n998 20.5561
R1405 VDPWR.n997 VDPWR.n966 20.5561
R1406 VDPWR.n1013 VDPWR.n1012 20.5561
R1407 VDPWR.n1016 VDPWR.n964 20.5561
R1408 VDPWR.n1017 VDPWR.n1016 20.5561
R1409 VDPWR.n1015 VDPWR.n962 20.5561
R1410 VDPWR.n1031 VDPWR.n1030 20.5561
R1411 VDPWR.n1034 VDPWR.n960 20.5561
R1412 VDPWR.n1035 VDPWR.n1034 20.5561
R1413 VDPWR.n1033 VDPWR.n958 20.5561
R1414 VDPWR.n1049 VDPWR.n1048 20.5561
R1415 VDPWR.n1052 VDPWR.n956 20.5561
R1416 VDPWR.n1053 VDPWR.n1052 20.5561
R1417 VDPWR.n1051 VDPWR.n954 20.5561
R1418 VDPWR.n1067 VDPWR.n1066 20.5561
R1419 VDPWR.n1070 VDPWR.n952 20.5561
R1420 VDPWR.n1071 VDPWR.n1070 20.5561
R1421 VDPWR.n1069 VDPWR.n950 20.5561
R1422 VDPWR.n1085 VDPWR.n1084 20.5561
R1423 VDPWR.n1088 VDPWR.n948 20.5561
R1424 VDPWR.n1089 VDPWR.n1088 20.5561
R1425 VDPWR.n1087 VDPWR.n946 20.5561
R1426 VDPWR.n1103 VDPWR.n1102 20.5561
R1427 VDPWR.n1106 VDPWR.n944 20.5561
R1428 VDPWR.n1107 VDPWR.n1106 20.5561
R1429 VDPWR.n1105 VDPWR.n942 20.5561
R1430 VDPWR.n833 VDPWR.n774 20.5561
R1431 VDPWR.n839 VDPWR.n833 20.5561
R1432 VDPWR.n831 VDPWR.n771 20.5561
R1433 VDPWR.n839 VDPWR.n831 20.5561
R1434 VDPWR.n829 VDPWR.n767 20.5561
R1435 VDPWR.n839 VDPWR.n829 20.5561
R1436 VDPWR.n827 VDPWR.n764 20.5561
R1437 VDPWR.n839 VDPWR.n827 20.5561
R1438 VDPWR.n825 VDPWR.n760 20.5561
R1439 VDPWR.n839 VDPWR.n825 20.5561
R1440 VDPWR.n823 VDPWR.n757 20.5561
R1441 VDPWR.n839 VDPWR.n823 20.5561
R1442 VDPWR.n821 VDPWR.n753 20.5561
R1443 VDPWR.n839 VDPWR.n821 20.5561
R1444 VDPWR.n819 VDPWR.n750 20.5561
R1445 VDPWR.n839 VDPWR.n819 20.5561
R1446 VDPWR.n817 VDPWR.n746 20.5561
R1447 VDPWR.n839 VDPWR.n817 20.5561
R1448 VDPWR.n815 VDPWR.n743 20.5561
R1449 VDPWR.n839 VDPWR.n815 20.5561
R1450 VDPWR.n813 VDPWR.n739 20.5561
R1451 VDPWR.n839 VDPWR.n813 20.5561
R1452 VDPWR.n811 VDPWR.n736 20.5561
R1453 VDPWR.n839 VDPWR.n811 20.5561
R1454 VDPWR.n809 VDPWR.n732 20.5561
R1455 VDPWR.n839 VDPWR.n809 20.5561
R1456 VDPWR.n807 VDPWR.n729 20.5561
R1457 VDPWR.n839 VDPWR.n807 20.5561
R1458 VDPWR.n805 VDPWR.n725 20.5561
R1459 VDPWR.n839 VDPWR.n805 20.5561
R1460 VDPWR.n803 VDPWR.n722 20.5561
R1461 VDPWR.n839 VDPWR.n803 20.5561
R1462 VDPWR.n801 VDPWR.n718 20.5561
R1463 VDPWR.n839 VDPWR.n801 20.5561
R1464 VDPWR.n799 VDPWR.n715 20.5561
R1465 VDPWR.n839 VDPWR.n799 20.5561
R1466 VDPWR.n797 VDPWR.n711 20.5561
R1467 VDPWR.n839 VDPWR.n797 20.5561
R1468 VDPWR.n795 VDPWR.n708 20.5561
R1469 VDPWR.n839 VDPWR.n795 20.5561
R1470 VDPWR.n793 VDPWR.n704 20.5561
R1471 VDPWR.n839 VDPWR.n793 20.5561
R1472 VDPWR.n791 VDPWR.n701 20.5561
R1473 VDPWR.n839 VDPWR.n791 20.5561
R1474 VDPWR.n789 VDPWR.n697 20.5561
R1475 VDPWR.n839 VDPWR.n789 20.5561
R1476 VDPWR.n787 VDPWR.n694 20.5561
R1477 VDPWR.n839 VDPWR.n787 20.5561
R1478 VDPWR.n785 VDPWR.n690 20.5561
R1479 VDPWR.n839 VDPWR.n785 20.5561
R1480 VDPWR.n783 VDPWR.n687 20.5561
R1481 VDPWR.n839 VDPWR.n783 20.5561
R1482 VDPWR.n838 VDPWR.n778 20.5561
R1483 VDPWR.n839 VDPWR.n838 20.5561
R1484 VDPWR.n835 VDPWR.n781 20.5561
R1485 VDPWR.n839 VDPWR.n835 20.5561
R1486 VDPWR.n841 VDPWR.n840 20.5561
R1487 VDPWR.n840 VDPWR.n839 20.5561
R1488 VDPWR.n492 VDPWR.n491 20.5561
R1489 VDPWR.n493 VDPWR.n492 20.5561
R1490 VDPWR.n180 VDPWR.n179 20.5561
R1491 VDPWR.n493 VDPWR.n180 20.5561
R1492 VDPWR.n503 VDPWR.n502 20.5561
R1493 VDPWR.n504 VDPWR.n503 20.5561
R1494 VDPWR.n174 VDPWR.n173 20.5561
R1495 VDPWR.n504 VDPWR.n174 20.5561
R1496 VDPWR.n190 VDPWR.n188 20.5561
R1497 VDPWR.n188 VDPWR.n186 20.5561
R1498 VDPWR.n189 VDPWR.n187 20.5561
R1499 VDPWR.n187 VDPWR.n186 20.5561
R1500 VDPWR.n184 VDPWR.n183 20.5561
R1501 VDPWR.n186 VDPWR.n184 20.5561
R1502 VDPWR.n185 VDPWR.n181 20.5561
R1503 VDPWR.n186 VDPWR.n185 20.5561
R1504 VDPWR.n214 VDPWR.n212 20.5561
R1505 VDPWR.n212 VDPWR.n210 20.5561
R1506 VDPWR.n213 VDPWR.n211 20.5561
R1507 VDPWR.n211 VDPWR.n210 20.5561
R1508 VDPWR.n208 VDPWR.n207 20.5561
R1509 VDPWR.n210 VDPWR.n208 20.5561
R1510 VDPWR.n209 VDPWR.n205 20.5561
R1511 VDPWR.n210 VDPWR.n209 20.5561
R1512 VDPWR.n238 VDPWR.n236 20.5561
R1513 VDPWR.n236 VDPWR.n234 20.5561
R1514 VDPWR.n237 VDPWR.n235 20.5561
R1515 VDPWR.n235 VDPWR.n234 20.5561
R1516 VDPWR.n232 VDPWR.n231 20.5561
R1517 VDPWR.n234 VDPWR.n232 20.5561
R1518 VDPWR.n233 VDPWR.n229 20.5561
R1519 VDPWR.n234 VDPWR.n233 20.5561
R1520 VDPWR.n262 VDPWR.n260 20.5561
R1521 VDPWR.n260 VDPWR.n258 20.5561
R1522 VDPWR.n261 VDPWR.n259 20.5561
R1523 VDPWR.n259 VDPWR.n258 20.5561
R1524 VDPWR.n256 VDPWR.n255 20.5561
R1525 VDPWR.n258 VDPWR.n256 20.5561
R1526 VDPWR.n257 VDPWR.n253 20.5561
R1527 VDPWR.n258 VDPWR.n257 20.5561
R1528 VDPWR.n286 VDPWR.n284 20.5561
R1529 VDPWR.n284 VDPWR.n282 20.5561
R1530 VDPWR.n285 VDPWR.n283 20.5561
R1531 VDPWR.n283 VDPWR.n282 20.5561
R1532 VDPWR.n280 VDPWR.n279 20.5561
R1533 VDPWR.n282 VDPWR.n280 20.5561
R1534 VDPWR.n281 VDPWR.n277 20.5561
R1535 VDPWR.n282 VDPWR.n281 20.5561
R1536 VDPWR.n310 VDPWR.n308 20.5561
R1537 VDPWR.n308 VDPWR.n306 20.5561
R1538 VDPWR.n309 VDPWR.n307 20.5561
R1539 VDPWR.n307 VDPWR.n306 20.5561
R1540 VDPWR.n304 VDPWR.n303 20.5561
R1541 VDPWR.n306 VDPWR.n304 20.5561
R1542 VDPWR.n305 VDPWR.n301 20.5561
R1543 VDPWR.n306 VDPWR.n305 20.5561
R1544 VDPWR.n154 VDPWR.n151 20.5561
R1545 VDPWR.n155 VDPWR.n154 20.5561
R1546 VDPWR.n131 VDPWR.n130 20.5561
R1547 VDPWR.n132 VDPWR.n131 20.5561
R1548 VDPWR.n11 VDPWR.n10 20.5561
R1549 VDPWR.n132 VDPWR.n11 20.5561
R1550 VDPWR.n142 VDPWR.n141 20.5561
R1551 VDPWR.n143 VDPWR.n142 20.5561
R1552 VDPWR.n5 VDPWR.n4 20.5561
R1553 VDPWR.n143 VDPWR.n5 20.5561
R1554 VDPWR.n21 VDPWR.n19 20.5561
R1555 VDPWR.n19 VDPWR.n17 20.5561
R1556 VDPWR.n20 VDPWR.n18 20.5561
R1557 VDPWR.n18 VDPWR.n17 20.5561
R1558 VDPWR.n15 VDPWR.n14 20.5561
R1559 VDPWR.n17 VDPWR.n15 20.5561
R1560 VDPWR.n16 VDPWR.n12 20.5561
R1561 VDPWR.n17 VDPWR.n16 20.5561
R1562 VDPWR.n40 VDPWR.n36 20.5561
R1563 VDPWR.n41 VDPWR.n40 20.5561
R1564 VDPWR.n39 VDPWR.n38 20.5561
R1565 VDPWR.n41 VDPWR.n39 20.5561
R1566 VDPWR.n45 VDPWR.n43 20.5561
R1567 VDPWR.n43 VDPWR.n41 20.5561
R1568 VDPWR.n44 VDPWR.n42 20.5561
R1569 VDPWR.n42 VDPWR.n41 20.5561
R1570 VDPWR.n1550 VDPWR.n1549 20.5561
R1571 VDPWR.n1549 VDPWR.n1548 20.5561
R1572 VDPWR.n1538 VDPWR.n1537 19.3338
R1573 VDPWR.n1537 VDPWR.n1536 19.3338
R1574 VDPWR.n1536 VDPWR.n1471 19.3338
R1575 VDPWR.n1531 VDPWR.n1471 19.3338
R1576 VDPWR.n1531 VDPWR.n1530 19.3338
R1577 VDPWR.n1530 VDPWR.n1529 19.3338
R1578 VDPWR.n1529 VDPWR.n1478 19.3338
R1579 VDPWR.n1524 VDPWR.n1478 19.3338
R1580 VDPWR.n1524 VDPWR.n1523 19.3338
R1581 VDPWR.n1523 VDPWR.n1522 19.3338
R1582 VDPWR.n1522 VDPWR.n1485 19.3338
R1583 VDPWR.n1506 VDPWR.n1485 19.3338
R1584 VDPWR.n1513 VDPWR.n1506 19.3338
R1585 VDPWR.n1513 VDPWR.n1512 19.3338
R1586 VDPWR.n939 VDPWR.n938 19.3338
R1587 VDPWR.n938 VDPWR.n937 19.3338
R1588 VDPWR.n937 VDPWR.n692 19.3338
R1589 VDPWR.n932 VDPWR.n692 19.3338
R1590 VDPWR.n932 VDPWR.n931 19.3338
R1591 VDPWR.n931 VDPWR.n930 19.3338
R1592 VDPWR.n930 VDPWR.n699 19.3338
R1593 VDPWR.n925 VDPWR.n699 19.3338
R1594 VDPWR.n925 VDPWR.n924 19.3338
R1595 VDPWR.n924 VDPWR.n923 19.3338
R1596 VDPWR.n923 VDPWR.n706 19.3338
R1597 VDPWR.n918 VDPWR.n706 19.3338
R1598 VDPWR.n918 VDPWR.n917 19.3338
R1599 VDPWR.n917 VDPWR.n916 19.3338
R1600 VDPWR.n916 VDPWR.n713 19.3338
R1601 VDPWR.n911 VDPWR.n713 19.3338
R1602 VDPWR.n911 VDPWR.n910 19.3338
R1603 VDPWR.n910 VDPWR.n909 19.3338
R1604 VDPWR.n909 VDPWR.n720 19.3338
R1605 VDPWR.n904 VDPWR.n720 19.3338
R1606 VDPWR.n904 VDPWR.n903 19.3338
R1607 VDPWR.n903 VDPWR.n902 19.3338
R1608 VDPWR.n902 VDPWR.n727 19.3338
R1609 VDPWR.n897 VDPWR.n727 19.3338
R1610 VDPWR.n897 VDPWR.n896 19.3338
R1611 VDPWR.n896 VDPWR.n895 19.3338
R1612 VDPWR.n895 VDPWR.n734 19.3338
R1613 VDPWR.n890 VDPWR.n734 19.3338
R1614 VDPWR.n890 VDPWR.n889 19.3338
R1615 VDPWR.n889 VDPWR.n888 19.3338
R1616 VDPWR.n888 VDPWR.n741 19.3338
R1617 VDPWR.n883 VDPWR.n741 19.3338
R1618 VDPWR.n883 VDPWR.n882 19.3338
R1619 VDPWR.n882 VDPWR.n881 19.3338
R1620 VDPWR.n881 VDPWR.n748 19.3338
R1621 VDPWR.n876 VDPWR.n748 19.3338
R1622 VDPWR.n876 VDPWR.n875 19.3338
R1623 VDPWR.n875 VDPWR.n874 19.3338
R1624 VDPWR.n874 VDPWR.n755 19.3338
R1625 VDPWR.n869 VDPWR.n755 19.3338
R1626 VDPWR.n869 VDPWR.n868 19.3338
R1627 VDPWR.n868 VDPWR.n867 19.3338
R1628 VDPWR.n867 VDPWR.n762 19.3338
R1629 VDPWR.n862 VDPWR.n762 19.3338
R1630 VDPWR.n862 VDPWR.n861 19.3338
R1631 VDPWR.n861 VDPWR.n860 19.3338
R1632 VDPWR.n860 VDPWR.n769 19.3338
R1633 VDPWR.n855 VDPWR.n769 19.3338
R1634 VDPWR.n855 VDPWR.n854 19.3338
R1635 VDPWR.n854 VDPWR.n853 19.3338
R1636 VDPWR.n853 VDPWR.n776 19.3338
R1637 VDPWR.n848 VDPWR.n776 19.3338
R1638 VDPWR.n848 VDPWR.n847 19.3338
R1639 VDPWR.n847 VDPWR.n846 19.3338
R1640 VDPWR.n678 VDPWR.n676 18.5005
R1641 VDPWR.n682 VDPWR.n676 18.5005
R1642 VDPWR.n661 VDPWR.n659 18.5005
R1643 VDPWR.n665 VDPWR.n659 18.5005
R1644 VDPWR.n644 VDPWR.n642 18.5005
R1645 VDPWR.n648 VDPWR.n642 18.5005
R1646 VDPWR.n627 VDPWR.n625 18.5005
R1647 VDPWR.n631 VDPWR.n625 18.5005
R1648 VDPWR.n610 VDPWR.n608 18.5005
R1649 VDPWR.n614 VDPWR.n608 18.5005
R1650 VDPWR.n593 VDPWR.n591 18.5005
R1651 VDPWR.n597 VDPWR.n591 18.5005
R1652 VDPWR.n576 VDPWR.n574 18.5005
R1653 VDPWR.n580 VDPWR.n574 18.5005
R1654 VDPWR.n559 VDPWR.n557 18.5005
R1655 VDPWR.n563 VDPWR.n557 18.5005
R1656 VDPWR.n565 VDPWR.n564 18.5005
R1657 VDPWR.n564 VDPWR.n563 18.5005
R1658 VDPWR.n582 VDPWR.n581 18.5005
R1659 VDPWR.n581 VDPWR.n580 18.5005
R1660 VDPWR.n599 VDPWR.n598 18.5005
R1661 VDPWR.n598 VDPWR.n597 18.5005
R1662 VDPWR.n616 VDPWR.n615 18.5005
R1663 VDPWR.n615 VDPWR.n614 18.5005
R1664 VDPWR.n633 VDPWR.n632 18.5005
R1665 VDPWR.n632 VDPWR.n631 18.5005
R1666 VDPWR.n650 VDPWR.n649 18.5005
R1667 VDPWR.n649 VDPWR.n648 18.5005
R1668 VDPWR.n667 VDPWR.n666 18.5005
R1669 VDPWR.n666 VDPWR.n665 18.5005
R1670 VDPWR.n684 VDPWR.n683 18.5005
R1671 VDPWR.n683 VDPWR.n682 18.5005
R1672 VDPWR.n467 VDPWR.n466 18.5005
R1673 VDPWR.n468 VDPWR.n467 18.5005
R1674 VDPWR.n202 VDPWR.n201 18.5005
R1675 VDPWR.n196 VDPWR.n195 18.5005
R1676 VDPWR.n469 VDPWR.n196 18.5005
R1677 VDPWR.n197 VDPWR.n191 18.5005
R1678 VDPWR.n441 VDPWR.n440 18.5005
R1679 VDPWR.n442 VDPWR.n441 18.5005
R1680 VDPWR.n226 VDPWR.n225 18.5005
R1681 VDPWR.n220 VDPWR.n219 18.5005
R1682 VDPWR.n443 VDPWR.n220 18.5005
R1683 VDPWR.n221 VDPWR.n215 18.5005
R1684 VDPWR.n415 VDPWR.n414 18.5005
R1685 VDPWR.n416 VDPWR.n415 18.5005
R1686 VDPWR.n250 VDPWR.n249 18.5005
R1687 VDPWR.n244 VDPWR.n243 18.5005
R1688 VDPWR.n417 VDPWR.n244 18.5005
R1689 VDPWR.n245 VDPWR.n239 18.5005
R1690 VDPWR.n389 VDPWR.n388 18.5005
R1691 VDPWR.n390 VDPWR.n389 18.5005
R1692 VDPWR.n274 VDPWR.n273 18.5005
R1693 VDPWR.n268 VDPWR.n267 18.5005
R1694 VDPWR.n391 VDPWR.n268 18.5005
R1695 VDPWR.n269 VDPWR.n263 18.5005
R1696 VDPWR.n363 VDPWR.n362 18.5005
R1697 VDPWR.n364 VDPWR.n363 18.5005
R1698 VDPWR.n298 VDPWR.n297 18.5005
R1699 VDPWR.n292 VDPWR.n291 18.5005
R1700 VDPWR.n365 VDPWR.n292 18.5005
R1701 VDPWR.n293 VDPWR.n287 18.5005
R1702 VDPWR.n329 VDPWR.n328 18.5005
R1703 VDPWR.n330 VDPWR.n329 18.5005
R1704 VDPWR.n322 VDPWR.n321 18.5005
R1705 VDPWR.n316 VDPWR.n315 18.5005
R1706 VDPWR.n331 VDPWR.n316 18.5005
R1707 VDPWR.n317 VDPWR.n311 18.5005
R1708 VDPWR.n98 VDPWR.n97 18.5005
R1709 VDPWR.n99 VDPWR.n98 18.5005
R1710 VDPWR.n33 VDPWR.n32 18.5005
R1711 VDPWR.n27 VDPWR.n26 18.5005
R1712 VDPWR.n100 VDPWR.n27 18.5005
R1713 VDPWR.n28 VDPWR.n22 18.5005
R1714 VDPWR.n64 VDPWR.n63 18.5005
R1715 VDPWR.n65 VDPWR.n64 18.5005
R1716 VDPWR.n57 VDPWR.n56 18.5005
R1717 VDPWR.n51 VDPWR.n50 18.5005
R1718 VDPWR.n66 VDPWR.n51 18.5005
R1719 VDPWR.n52 VDPWR.n46 18.5005
R1720 VDPWR.n164 VDPWR.n163 18.5005
R1721 VDPWR.n1170 VDPWR.n1169 16.8187
R1722 VDPWR.n1172 VDPWR.n1171 16.8187
R1723 VDPWR.n1166 VDPWR.n1159 16.8187
R1724 VDPWR.n1173 VDPWR.n1166 16.8187
R1725 VDPWR.n1186 VDPWR.n1184 16.8187
R1726 VDPWR.n1187 VDPWR.n1154 16.8187
R1727 VDPWR.n1188 VDPWR.n1187 16.8187
R1728 VDPWR.n1202 VDPWR.n1200 16.8187
R1729 VDPWR.n1203 VDPWR.n1149 16.8187
R1730 VDPWR.n1204 VDPWR.n1203 16.8187
R1731 VDPWR.n1218 VDPWR.n1216 16.8187
R1732 VDPWR.n1219 VDPWR.n1144 16.8187
R1733 VDPWR.n1220 VDPWR.n1219 16.8187
R1734 VDPWR.n1234 VDPWR.n1232 16.8187
R1735 VDPWR.n1235 VDPWR.n1139 16.8187
R1736 VDPWR.n1236 VDPWR.n1235 16.8187
R1737 VDPWR.n1250 VDPWR.n1248 16.8187
R1738 VDPWR.n1251 VDPWR.n1134 16.8187
R1739 VDPWR.n1252 VDPWR.n1251 16.8187
R1740 VDPWR.n1266 VDPWR.n1264 16.8187
R1741 VDPWR.n1267 VDPWR.n1129 16.8187
R1742 VDPWR.n1268 VDPWR.n1267 16.8187
R1743 VDPWR.n1282 VDPWR.n1280 16.8187
R1744 VDPWR.n1283 VDPWR.n1124 16.8187
R1745 VDPWR.n1284 VDPWR.n1283 16.8187
R1746 VDPWR.n1298 VDPWR.n1296 16.8187
R1747 VDPWR.n1299 VDPWR.n1119 16.8187
R1748 VDPWR.n1300 VDPWR.n1299 16.8187
R1749 VDPWR.n566 VDPWR.n551 16.8187
R1750 VDPWR.n554 VDPWR.n551 16.8187
R1751 VDPWR.n583 VDPWR.n546 16.8187
R1752 VDPWR.n571 VDPWR.n546 16.8187
R1753 VDPWR.n600 VDPWR.n541 16.8187
R1754 VDPWR.n588 VDPWR.n541 16.8187
R1755 VDPWR.n617 VDPWR.n536 16.8187
R1756 VDPWR.n605 VDPWR.n536 16.8187
R1757 VDPWR.n634 VDPWR.n531 16.8187
R1758 VDPWR.n622 VDPWR.n531 16.8187
R1759 VDPWR.n651 VDPWR.n526 16.8187
R1760 VDPWR.n639 VDPWR.n526 16.8187
R1761 VDPWR.n668 VDPWR.n521 16.8187
R1762 VDPWR.n656 VDPWR.n521 16.8187
R1763 VDPWR.n685 VDPWR.n516 16.8187
R1764 VDPWR.n673 VDPWR.n516 16.8187
R1765 VDPWR.n1456 VDPWR.n1311 16.8187
R1766 VDPWR.n1457 VDPWR.n1456 16.8187
R1767 VDPWR.n1454 VDPWR.n1316 16.8187
R1768 VDPWR.n1455 VDPWR.n1454 16.8187
R1769 VDPWR.n1452 VDPWR.n1451 16.8187
R1770 VDPWR.n1453 VDPWR.n1452 16.8187
R1771 VDPWR.n1430 VDPWR.n1323 16.8187
R1772 VDPWR.n1431 VDPWR.n1430 16.8187
R1773 VDPWR.n1432 VDPWR.n1327 16.8187
R1774 VDPWR.n1433 VDPWR.n1432 16.8187
R1775 VDPWR.n1426 VDPWR.n1332 16.8187
R1776 VDPWR.n1427 VDPWR.n1426 16.8187
R1777 VDPWR.n1424 VDPWR.n1423 16.8187
R1778 VDPWR.n1425 VDPWR.n1424 16.8187
R1779 VDPWR.n1402 VDPWR.n1339 16.8187
R1780 VDPWR.n1403 VDPWR.n1402 16.8187
R1781 VDPWR.n1404 VDPWR.n1343 16.8187
R1782 VDPWR.n1405 VDPWR.n1404 16.8187
R1783 VDPWR.n1398 VDPWR.n1348 16.8187
R1784 VDPWR.n1399 VDPWR.n1398 16.8187
R1785 VDPWR.n1396 VDPWR.n1395 16.8187
R1786 VDPWR.n1397 VDPWR.n1396 16.8187
R1787 VDPWR.n1376 VDPWR.n1355 16.8187
R1788 VDPWR.n1377 VDPWR.n1376 16.8187
R1789 VDPWR.n1373 VDPWR.n1372 16.8187
R1790 VDPWR.n1366 VDPWR.n1359 16.8187
R1791 VDPWR.n1378 VDPWR.n1366 16.8187
R1792 VDPWR.n1371 VDPWR.n1370 16.8187
R1793 VDPWR.n565 VDPWR.n552 14.3397
R1794 VDPWR.n582 VDPWR.n569 14.3397
R1795 VDPWR.n599 VDPWR.n586 14.3397
R1796 VDPWR.n616 VDPWR.n603 14.3397
R1797 VDPWR.n633 VDPWR.n620 14.3397
R1798 VDPWR.n650 VDPWR.n637 14.3397
R1799 VDPWR.n667 VDPWR.n654 14.3397
R1800 VDPWR.n684 VDPWR.n671 14.3397
R1801 VDPWR.n680 VDPWR.n678 13.8537
R1802 VDPWR.n678 VDPWR.n671 13.8537
R1803 VDPWR.n663 VDPWR.n661 13.8537
R1804 VDPWR.n661 VDPWR.n654 13.8537
R1805 VDPWR.n646 VDPWR.n644 13.8537
R1806 VDPWR.n644 VDPWR.n637 13.8537
R1807 VDPWR.n629 VDPWR.n627 13.8537
R1808 VDPWR.n627 VDPWR.n620 13.8537
R1809 VDPWR.n612 VDPWR.n610 13.8537
R1810 VDPWR.n610 VDPWR.n603 13.8537
R1811 VDPWR.n595 VDPWR.n593 13.8537
R1812 VDPWR.n593 VDPWR.n586 13.8537
R1813 VDPWR.n578 VDPWR.n576 13.8537
R1814 VDPWR.n576 VDPWR.n569 13.8537
R1815 VDPWR.n561 VDPWR.n559 13.8537
R1816 VDPWR.n559 VDPWR.n552 13.8537
R1817 VDPWR.n679 VDPWR.n675 13.2148
R1818 VDPWR.n662 VDPWR.n658 13.2148
R1819 VDPWR.n645 VDPWR.n641 13.2148
R1820 VDPWR.n628 VDPWR.n624 13.2148
R1821 VDPWR.n611 VDPWR.n607 13.2148
R1822 VDPWR.n594 VDPWR.n590 13.2148
R1823 VDPWR.n577 VDPWR.n573 13.2148
R1824 VDPWR.n560 VDPWR.n556 13.2148
R1825 VDPWR.n511 VDPWR.n168 12.6054
R1826 VDPWR.n1176 VDPWR.n1175 11.563
R1827 VDPWR.n1175 VDPWR.n1174 11.563
R1828 VDPWR.n1189 VDPWR.n1185 11.563
R1829 VDPWR.n1205 VDPWR.n1201 11.563
R1830 VDPWR.n1221 VDPWR.n1217 11.563
R1831 VDPWR.n1237 VDPWR.n1233 11.563
R1832 VDPWR.n1253 VDPWR.n1249 11.563
R1833 VDPWR.n1269 VDPWR.n1265 11.563
R1834 VDPWR.n1285 VDPWR.n1281 11.563
R1835 VDPWR.n1301 VDPWR.n1297 11.563
R1836 VDPWR.n1458 VDPWR.n1317 11.563
R1837 VDPWR.n1428 VDPWR.n1318 11.563
R1838 VDPWR.n1434 VDPWR.n1333 11.563
R1839 VDPWR.n1400 VDPWR.n1334 11.563
R1840 VDPWR.n1406 VDPWR.n1349 11.563
R1841 VDPWR.n1374 VDPWR.n1350 11.563
R1842 VDPWR.n1381 VDPWR.n1380 11.563
R1843 VDPWR.n1380 VDPWR.n1379 11.563
R1844 VDPWR.n1191 VDPWR.n1185 10.2708
R1845 VDPWR.n1207 VDPWR.n1201 10.2708
R1846 VDPWR.n1223 VDPWR.n1217 10.2708
R1847 VDPWR.n1239 VDPWR.n1233 10.2708
R1848 VDPWR.n1255 VDPWR.n1249 10.2708
R1849 VDPWR.n1271 VDPWR.n1265 10.2708
R1850 VDPWR.n1287 VDPWR.n1281 10.2708
R1851 VDPWR.n1303 VDPWR.n1297 10.2708
R1852 VDPWR.n1460 VDPWR.n1317 10.2708
R1853 VDPWR.n1324 VDPWR.n1318 10.2708
R1854 VDPWR.n1436 VDPWR.n1333 10.2708
R1855 VDPWR.n1340 VDPWR.n1334 10.2708
R1856 VDPWR.n1408 VDPWR.n1349 10.2708
R1857 VDPWR.n1356 VDPWR.n1350 10.2708
R1858 VDPWR.n1362 VDPWR.t19 9.52217
R1859 VDPWR.n1362 VDPWR.t17 9.52217
R1860 VDPWR.n1361 VDPWR.t575 9.52217
R1861 VDPWR.n1361 VDPWR.t52 9.52217
R1862 VDPWR.n1360 VDPWR.t359 9.52217
R1863 VDPWR.n1360 VDPWR.t181 9.52217
R1864 VDPWR.n1358 VDPWR.t546 9.52217
R1865 VDPWR.n1358 VDPWR.t270 9.52217
R1866 VDPWR.n1357 VDPWR.t253 9.52217
R1867 VDPWR.n1357 VDPWR.t544 9.52217
R1868 VDPWR.n1389 VDPWR.t234 9.52217
R1869 VDPWR.n1389 VDPWR.t56 9.52217
R1870 VDPWR.n1390 VDPWR.t117 9.52217
R1871 VDPWR.n1390 VDPWR.t540 9.52217
R1872 VDPWR.n1351 VDPWR.t351 9.52217
R1873 VDPWR.n1351 VDPWR.t487 9.52217
R1874 VDPWR.n1346 VDPWR.t481 9.52217
R1875 VDPWR.n1346 VDPWR.t353 9.52217
R1876 VDPWR.n1345 VDPWR.t542 9.52217
R1877 VDPWR.n1345 VDPWR.t158 9.52217
R1878 VDPWR.n1344 VDPWR.t152 9.52217
R1879 VDPWR.n1344 VDPWR.t121 9.52217
R1880 VDPWR.n1342 VDPWR.t375 9.52217
R1881 VDPWR.n1342 VDPWR.t531 9.52217
R1882 VDPWR.n1341 VDPWR.t76 9.52217
R1883 VDPWR.n1341 VDPWR.t519 9.52217
R1884 VDPWR.n1417 VDPWR.t304 9.52217
R1885 VDPWR.n1417 VDPWR.t308 9.52217
R1886 VDPWR.n1418 VDPWR.t306 9.52217
R1887 VDPWR.n1418 VDPWR.t380 9.52217
R1888 VDPWR.n1335 VDPWR.t585 9.52217
R1889 VDPWR.n1335 VDPWR.t272 9.52217
R1890 VDPWR.n1330 VDPWR.t344 9.52217
R1891 VDPWR.n1330 VDPWR.t276 9.52217
R1892 VDPWR.n1329 VDPWR.t40 9.52217
R1893 VDPWR.n1329 VDPWR.t96 9.52217
R1894 VDPWR.n1328 VDPWR.t314 9.52217
R1895 VDPWR.n1328 VDPWR.t213 9.52217
R1896 VDPWR.n1326 VDPWR.t88 9.52217
R1897 VDPWR.n1326 VDPWR.t366 9.52217
R1898 VDPWR.n1325 VDPWR.t74 9.52217
R1899 VDPWR.n1325 VDPWR.t127 9.52217
R1900 VDPWR.n1445 VDPWR.t413 9.52217
R1901 VDPWR.n1445 VDPWR.t92 9.52217
R1902 VDPWR.n1446 VDPWR.t90 9.52217
R1903 VDPWR.n1446 VDPWR.t415 9.52217
R1904 VDPWR.n1319 VDPWR.t54 9.52217
R1905 VDPWR.n1319 VDPWR.t423 9.52217
R1906 VDPWR.n1314 VDPWR.t421 9.52217
R1907 VDPWR.n1314 VDPWR.t300 9.52217
R1908 VDPWR.n1313 VDPWR.t506 9.52217
R1909 VDPWR.n1313 VDPWR.t50 9.52217
R1910 VDPWR.n1312 VDPWR.t201 9.52217
R1911 VDPWR.n1312 VDPWR.t230 9.52217
R1912 VDPWR.n1167 VDPWR.t471 9.52217
R1913 VDPWR.n1167 VDPWR.t536 9.52217
R1914 VDPWR.n1162 VDPWR.t133 9.52217
R1915 VDPWR.n1162 VDPWR.t228 9.52217
R1916 VDPWR.n1161 VDPWR.t175 9.52217
R1917 VDPWR.n1161 VDPWR.t36 9.52217
R1918 VDPWR.n1160 VDPWR.t349 9.52217
R1919 VDPWR.n1160 VDPWR.t177 9.52217
R1920 VDPWR.n1181 VDPWR.t548 9.52217
R1921 VDPWR.n1181 VDPWR.t552 9.52217
R1922 VDPWR.n1157 VDPWR.t550 9.52217
R1923 VDPWR.n1157 VDPWR.t278 9.52217
R1924 VDPWR.n1156 VDPWR.t571 9.52217
R1925 VDPWR.n1156 VDPWR.t569 9.52217
R1926 VDPWR.n1155 VDPWR.t524 9.52217
R1927 VDPWR.n1155 VDPWR.t364 9.52217
R1928 VDPWR.n1197 VDPWR.t195 9.52217
R1929 VDPWR.n1197 VDPWR.t517 9.52217
R1930 VDPWR.n1152 VDPWR.t377 9.52217
R1931 VDPWR.n1152 VDPWR.t240 9.52217
R1932 VDPWR.n1151 VDPWR.t255 9.52217
R1933 VDPWR.n1151 VDPWR.t312 9.52217
R1934 VDPWR.n1150 VDPWR.t310 9.52217
R1935 VDPWR.n1150 VDPWR.t257 9.52217
R1936 VDPWR.n1213 VDPWR.t62 9.52217
R1937 VDPWR.n1213 VDPWR.t538 9.52217
R1938 VDPWR.n1147 VDPWR.t232 9.52217
R1939 VDPWR.n1147 VDPWR.t86 9.52217
R1940 VDPWR.n1146 VDPWR.t48 9.52217
R1941 VDPWR.n1146 VDPWR.t496 9.52217
R1942 VDPWR.n1145 VDPWR.t80 9.52217
R1943 VDPWR.n1145 VDPWR.t68 9.52217
R1944 VDPWR.n1229 VDPWR.t282 9.52217
R1945 VDPWR.n1229 VDPWR.t42 9.52217
R1946 VDPWR.n1142 VDPWR.t191 9.52217
R1947 VDPWR.n1142 VDPWR.t189 9.52217
R1948 VDPWR.n1141 VDPWR.t477 9.52217
R1949 VDPWR.n1141 VDPWR.t475 9.52217
R1950 VDPWR.n1140 VDPWR.t298 9.52217
R1951 VDPWR.n1140 VDPWR.t484 9.52217
R1952 VDPWR.n1245 VDPWR.t294 9.52217
R1953 VDPWR.n1245 VDPWR.t288 9.52217
R1954 VDPWR.n1137 VDPWR.t290 9.52217
R1955 VDPWR.n1137 VDPWR.t292 9.52217
R1956 VDPWR.n1136 VDPWR.t604 9.52217
R1957 VDPWR.n1136 VDPWR.t396 9.52217
R1958 VDPWR.n1135 VDPWR.t296 9.52217
R1959 VDPWR.n1135 VDPWR.t394 9.52217
R1960 VDPWR.n1261 VDPWR.t527 9.52217
R1961 VDPWR.n1261 VDPWR.t119 9.52217
R1962 VDPWR.n1132 VDPWR.t60 9.52217
R1963 VDPWR.n1132 VDPWR.t58 9.52217
R1964 VDPWR.n1131 VDPWR.t407 9.52217
R1965 VDPWR.n1131 VDPWR.t411 9.52217
R1966 VDPWR.n1130 VDPWR.t431 9.52217
R1967 VDPWR.n1130 VDPWR.t409 9.52217
R1968 VDPWR.n1277 VDPWR.t109 9.52217
R1969 VDPWR.n1277 VDPWR.t38 9.52217
R1970 VDPWR.n1127 VDPWR.t429 9.52217
R1971 VDPWR.n1127 VDPWR.t107 9.52217
R1972 VDPWR.n1126 VDPWR.t46 9.52217
R1973 VDPWR.n1126 VDPWR.t529 9.52217
R1974 VDPWR.n1125 VDPWR.t614 9.52217
R1975 VDPWR.n1125 VDPWR.t44 9.52217
R1976 VDPWR.n1293 VDPWR.t13 9.52217
R1977 VDPWR.n1293 VDPWR.t564 9.52217
R1978 VDPWR.n1122 VDPWR.t11 9.52217
R1979 VDPWR.n1122 VDPWR.t5 9.52217
R1980 VDPWR.n1121 VDPWR.t342 9.52217
R1981 VDPWR.n1121 VDPWR.t268 9.52217
R1982 VDPWR.n1120 VDPWR.t66 9.52217
R1983 VDPWR.n1120 VDPWR.t225 9.52217
R1984 VDPWR.n974 VDPWR.t385 9.52217
R1985 VDPWR.n974 VDPWR.t170 9.52217
R1986 VDPWR.n971 VDPWR.t498 9.52217
R1987 VDPWR.n971 VDPWR.t578 9.52217
R1988 VDPWR.n991 VDPWR.t64 9.52217
R1989 VDPWR.n991 VDPWR.t370 9.52217
R1990 VDPWR.n967 VDPWR.t581 9.52217
R1991 VDPWR.n967 VDPWR.t168 9.52217
R1992 VDPWR.n1009 VDPWR.t398 9.52217
R1993 VDPWR.n1009 VDPWR.t115 9.52217
R1994 VDPWR.n963 VDPWR.t400 9.52217
R1995 VDPWR.n963 VDPWR.t249 9.52217
R1996 VDPWR.n1027 VDPWR.t146 9.52217
R1997 VDPWR.n1027 VDPWR.t236 9.52217
R1998 VDPWR.n959 VDPWR.t357 9.52217
R1999 VDPWR.n959 VDPWR.t238 9.52217
R2000 VDPWR.n1045 VDPWR.t185 9.52217
R2001 VDPWR.n1045 VDPWR.t362 9.52217
R2002 VDPWR.n955 VDPWR.t183 9.52217
R2003 VDPWR.n955 VDPWR.t156 9.52217
R2004 VDPWR.n1063 VDPWR.t320 9.52217
R2005 VDPWR.n1063 VDPWR.t323 9.52217
R2006 VDPWR.n951 VDPWR.t318 9.52217
R2007 VDPWR.n951 VDPWR.t325 9.52217
R2008 VDPWR.n1081 VDPWR.t203 9.52217
R2009 VDPWR.n1081 VDPWR.t425 9.52217
R2010 VDPWR.n947 VDPWR.t205 9.52217
R2011 VDPWR.n947 VDPWR.t587 9.52217
R2012 VDPWR.n1099 VDPWR.t274 9.52217
R2013 VDPWR.n1099 VDPWR.t70 9.52217
R2014 VDPWR.n943 VDPWR.t346 9.52217
R2015 VDPWR.n943 VDPWR.t600 9.52217
R2016 VDPWR.n1367 VDPWR.t15 9.52217
R2017 VDPWR.n1367 VDPWR.t94 9.52217
R2018 VDPWR.n203 VDPWR.t355 9.52217
R2019 VDPWR.n203 VDPWR.t419 9.52217
R2020 VDPWR.n192 VDPWR.t328 9.52217
R2021 VDPWR.n192 VDPWR.t562 9.52217
R2022 VDPWR.n227 VDPWR.t166 9.52217
R2023 VDPWR.n227 VDPWR.t135 9.52217
R2024 VDPWR.n216 VDPWR.t508 9.52217
R2025 VDPWR.n216 VDPWR.t131 9.52217
R2026 VDPWR.n251 VDPWR.t591 9.52217
R2027 VDPWR.n251 VDPWR.t338 9.52217
R2028 VDPWR.n240 VDPWR.t244 9.52217
R2029 VDPWR.n240 VDPWR.t242 9.52217
R2030 VDPWR.n275 VDPWR.t417 9.52217
R2031 VDPWR.n275 VDPWR.t286 9.52217
R2032 VDPWR.n264 VDPWR.t515 9.52217
R2033 VDPWR.n264 VDPWR.t336 9.52217
R2034 VDPWR.n299 VDPWR.t98 9.52217
R2035 VDPWR.n299 VDPWR.t30 9.52217
R2036 VDPWR.n288 VDPWR.t207 9.52217
R2037 VDPWR.n288 VDPWR.t221 9.52217
R2038 VDPWR.n323 VDPWR.t437 9.52217
R2039 VDPWR.n323 VDPWR.t449 9.52217
R2040 VDPWR.n312 VDPWR.t513 9.52217
R2041 VDPWR.n312 VDPWR.t149 9.52217
R2042 VDPWR.n34 VDPWR.t464 9.52217
R2043 VDPWR.n34 VDPWR.t440 9.52217
R2044 VDPWR.n23 VDPWR.t373 9.52217
R2045 VDPWR.n23 VDPWR.t23 9.52217
R2046 VDPWR.n58 VDPWR.t434 9.52217
R2047 VDPWR.n58 VDPWR.t446 9.52217
R2048 VDPWR.n47 VDPWR.t504 9.52217
R2049 VDPWR.n47 VDPWR.t502 9.52217
R2050 VDPWR.n1516 VDPWR.t82 9.39094
R2051 VDPWR.n156 VDPWR.n155 8.66346
R2052 VDPWR.n496 VDPWR.n495 7.70883
R2053 VDPWR.n507 VDPWR.n506 7.70883
R2054 VDPWR.n135 VDPWR.n134 7.70883
R2055 VDPWR.n146 VDPWR.n145 7.70883
R2056 VDPWR.n1548 VDPWR.n1547 7.4066
R2057 VDPWR.n496 VDPWR.n177 6.57828
R2058 VDPWR.n507 VDPWR.n171 6.57828
R2059 VDPWR.n135 VDPWR.n8 6.57828
R2060 VDPWR.n146 VDPWR.n2 6.57828
R2061 VDPWR.n985 VDPWR.n983 5.44168
R2062 VDPWR.n983 VDPWR.n982 5.44168
R2063 VDPWR.n1003 VDPWR.n1001 5.44168
R2064 VDPWR.n1001 VDPWR.n1000 5.44168
R2065 VDPWR.n1021 VDPWR.n1019 5.44168
R2066 VDPWR.n1019 VDPWR.n1018 5.44168
R2067 VDPWR.n1039 VDPWR.n1037 5.44168
R2068 VDPWR.n1037 VDPWR.n1036 5.44168
R2069 VDPWR.n1057 VDPWR.n1055 5.44168
R2070 VDPWR.n1055 VDPWR.n1054 5.44168
R2071 VDPWR.n1075 VDPWR.n1073 5.44168
R2072 VDPWR.n1073 VDPWR.n1072 5.44168
R2073 VDPWR.n1093 VDPWR.n1091 5.44168
R2074 VDPWR.n1091 VDPWR.n1090 5.44168
R2075 VDPWR.n1111 VDPWR.n1109 5.44168
R2076 VDPWR.n1109 VDPWR.n1108 5.44168
R2077 VDPWR.n494 VDPWR.n493 5.33119
R2078 VDPWR.n133 VDPWR.n132 5.33119
R2079 VDPWR.n505 VDPWR.n504 5.31424
R2080 VDPWR.n144 VDPWR.n143 5.31424
R2081 VDPWR.n1175 VDPWR.n1165 5.0005
R2082 VDPWR.n1380 VDPWR.n1365 5.0005
R2083 VDPWR.n1542 VDPWR.n1310 4.63898
R2084 VDPWR.n556 VDPWR.n555 4.40526
R2085 VDPWR.n573 VDPWR.n572 4.40526
R2086 VDPWR.n590 VDPWR.n589 4.40526
R2087 VDPWR.n607 VDPWR.n606 4.40526
R2088 VDPWR.n624 VDPWR.n623 4.40526
R2089 VDPWR.n641 VDPWR.n640 4.40526
R2090 VDPWR.n658 VDPWR.n657 4.40526
R2091 VDPWR.n675 VDPWR.n674 4.40526
R2092 VDPWR.n1542 VDPWR.n1541 4.29701
R2093 VDPWR.n1174 VDPWR.n1172 3.72599
R2094 VDPWR.n1190 VDPWR.n1189 3.72599
R2095 VDPWR.n1206 VDPWR.n1205 3.72599
R2096 VDPWR.n1222 VDPWR.n1221 3.72599
R2097 VDPWR.n1238 VDPWR.n1237 3.72599
R2098 VDPWR.n1254 VDPWR.n1253 3.72599
R2099 VDPWR.n1270 VDPWR.n1269 3.72599
R2100 VDPWR.n1286 VDPWR.n1285 3.72599
R2101 VDPWR.n1302 VDPWR.n1301 3.72599
R2102 VDPWR.n1379 VDPWR.n1373 3.72599
R2103 VDPWR.n1375 VDPWR.n1374 3.72599
R2104 VDPWR.n1407 VDPWR.n1406 3.72599
R2105 VDPWR.n1401 VDPWR.n1400 3.72599
R2106 VDPWR.n1435 VDPWR.n1434 3.72599
R2107 VDPWR.n1429 VDPWR.n1428 3.72599
R2108 VDPWR.n1459 VDPWR.n1458 3.72599
R2109 VDPWR.n1544 VDPWR.n511 3.30858
R2110 VDPWR.n1544 VDPWR.n1543 3.19848
R2111 VDPWR.n355 VDPWR.n354 3.13979
R2112 VDPWR.n124 VDPWR.n123 3.13979
R2113 VDPWR.n90 VDPWR.n89 3.13979
R2114 VDPWR.n1117 VDPWR 2.86795
R2115 VDPWR.n839 VDPWR.t24 2.77153
R2116 VDPWR.n976 VDPWR.n975 2.53478
R2117 VDPWR.n983 VDPWR.n978 2.35344
R2118 VDPWR.n1001 VDPWR.n996 2.35344
R2119 VDPWR.n1019 VDPWR.n1014 2.35344
R2120 VDPWR.n1037 VDPWR.n1032 2.35344
R2121 VDPWR.n1055 VDPWR.n1050 2.35344
R2122 VDPWR.n1073 VDPWR.n1068 2.35344
R2123 VDPWR.n1091 VDPWR.n1086 2.35344
R2124 VDPWR.n1109 VDPWR.n1104 2.35344
R2125 VDPWR.n1512 VDPWR.n1511 2.3255
R2126 VDPWR.n1506 VDPWR.n1487 2.3255
R2127 VDPWR.n846 VDPWR.n845 2.3255
R2128 VDPWR.n849 VDPWR.n848 2.3255
R2129 VDPWR.n853 VDPWR.n852 2.3255
R2130 VDPWR.n856 VDPWR.n855 2.3255
R2131 VDPWR.n860 VDPWR.n859 2.3255
R2132 VDPWR.n863 VDPWR.n862 2.3255
R2133 VDPWR.n867 VDPWR.n866 2.3255
R2134 VDPWR.n870 VDPWR.n869 2.3255
R2135 VDPWR.n874 VDPWR.n873 2.3255
R2136 VDPWR.n877 VDPWR.n876 2.3255
R2137 VDPWR.n881 VDPWR.n880 2.3255
R2138 VDPWR.n884 VDPWR.n883 2.3255
R2139 VDPWR.n888 VDPWR.n887 2.3255
R2140 VDPWR.n891 VDPWR.n890 2.3255
R2141 VDPWR.n895 VDPWR.n894 2.3255
R2142 VDPWR.n898 VDPWR.n897 2.3255
R2143 VDPWR.n902 VDPWR.n901 2.3255
R2144 VDPWR.n905 VDPWR.n904 2.3255
R2145 VDPWR.n909 VDPWR.n908 2.3255
R2146 VDPWR.n912 VDPWR.n911 2.3255
R2147 VDPWR.n916 VDPWR.n915 2.3255
R2148 VDPWR.n919 VDPWR.n918 2.3255
R2149 VDPWR.n923 VDPWR.n922 2.3255
R2150 VDPWR.n926 VDPWR.n925 2.3255
R2151 VDPWR.n930 VDPWR.n929 2.3255
R2152 VDPWR.n933 VDPWR.n932 2.3255
R2153 VDPWR.n937 VDPWR.n936 2.3255
R2154 VDPWR.n940 VDPWR.n939 2.3255
R2155 VDPWR.n1522 VDPWR.n1521 2.3255
R2156 VDPWR.n1525 VDPWR.n1524 2.3255
R2157 VDPWR.n1529 VDPWR.n1528 2.3255
R2158 VDPWR.n1532 VDPWR.n1531 2.3255
R2159 VDPWR.n1536 VDPWR.n1535 2.3255
R2160 VDPWR.n1539 VDPWR.n1538 2.3255
R2161 VDPWR.n347 VDPWR.n346 2.3255
R2162 VDPWR.n342 VDPWR.n341 2.3255
R2163 VDPWR.n381 VDPWR.n380 2.3255
R2164 VDPWR.n376 VDPWR.n375 2.3255
R2165 VDPWR.n407 VDPWR.n406 2.3255
R2166 VDPWR.n402 VDPWR.n401 2.3255
R2167 VDPWR.n433 VDPWR.n432 2.3255
R2168 VDPWR.n428 VDPWR.n427 2.3255
R2169 VDPWR.n459 VDPWR.n458 2.3255
R2170 VDPWR.n454 VDPWR.n453 2.3255
R2171 VDPWR.n485 VDPWR.n484 2.3255
R2172 VDPWR.n480 VDPWR.n479 2.3255
R2173 VDPWR.n159 VDPWR.n158 2.3255
R2174 VDPWR.n82 VDPWR.n81 2.3255
R2175 VDPWR.n77 VDPWR.n76 2.3255
R2176 VDPWR.n116 VDPWR.n115 2.3255
R2177 VDPWR.n111 VDPWR.n110 2.3255
R2178 VDPWR.n987 VDPWR.n972 2.29581
R2179 VDPWR.n990 VDPWR.n970 2.29581
R2180 VDPWR.n994 VDPWR.n993 2.29581
R2181 VDPWR.n1005 VDPWR.n968 2.29581
R2182 VDPWR.n1008 VDPWR.n966 2.29581
R2183 VDPWR.n1012 VDPWR.n1011 2.29581
R2184 VDPWR.n1023 VDPWR.n964 2.29581
R2185 VDPWR.n1026 VDPWR.n962 2.29581
R2186 VDPWR.n1030 VDPWR.n1029 2.29581
R2187 VDPWR.n1041 VDPWR.n960 2.29581
R2188 VDPWR.n1044 VDPWR.n958 2.29581
R2189 VDPWR.n1048 VDPWR.n1047 2.29581
R2190 VDPWR.n1059 VDPWR.n956 2.29581
R2191 VDPWR.n1062 VDPWR.n954 2.29581
R2192 VDPWR.n1066 VDPWR.n1065 2.29581
R2193 VDPWR.n1077 VDPWR.n952 2.29581
R2194 VDPWR.n1080 VDPWR.n950 2.29581
R2195 VDPWR.n1084 VDPWR.n1083 2.29581
R2196 VDPWR.n1095 VDPWR.n948 2.29581
R2197 VDPWR.n1098 VDPWR.n946 2.29581
R2198 VDPWR.n1102 VDPWR.n1101 2.29581
R2199 VDPWR.n1113 VDPWR.n944 2.29581
R2200 VDPWR.n1116 VDPWR.n942 2.29581
R2201 VDPWR.n357 VDPWR.n356 2.2505
R2202 VDPWR.n92 VDPWR.n91 2.2505
R2203 VDPWR.n126 VDPWR.n125 2.2505
R2204 VDPWR.n160 VDPWR.n151 2.2281
R2205 VDPWR.n1169 VDPWR.n1168 2.1858
R2206 VDPWR.n157 VDPWR.n152 2.17472
R2207 VDPWR.n1551 VDPWR.n1550 2.17342
R2208 VDPWR.n1546 VDPWR.n1545 2.17342
R2209 VDPWR.n1509 VDPWR.n1508 2.16821
R2210 VDPWR.n1514 VDPWR.n1504 2.16821
R2211 VDPWR.n1519 VDPWR.n1518 2.16821
R2212 VDPWR.n73 VDPWR.n44 2.16821
R2213 VDPWR.n567 VDPWR.n566 2.122
R2214 VDPWR.n584 VDPWR.n583 2.122
R2215 VDPWR.n601 VDPWR.n600 2.122
R2216 VDPWR.n618 VDPWR.n617 2.122
R2217 VDPWR.n635 VDPWR.n634 2.122
R2218 VDPWR.n652 VDPWR.n651 2.122
R2219 VDPWR.n669 VDPWR.n668 2.122
R2220 VDPWR.n686 VDPWR.n685 2.122
R2221 VDPWR.t20 VDPWR.t222 2.08383
R2222 VDPWR.t572 VDPWR.t77 2.08383
R2223 VDPWR.t0 VDPWR.t178 2.07474
R2224 VDPWR.t26 VDPWR.t472 2.07474
R2225 VDPWR.n1370 VDPWR.n1369 2.0647
R2226 VDPWR.n1540 VDPWR.n1466 2.04321
R2227 VDPWR.n1472 VDPWR.n1469 2.04321
R2228 VDPWR.n1533 VDPWR.n1473 2.04321
R2229 VDPWR.n1479 VDPWR.n1476 2.04321
R2230 VDPWR.n1526 VDPWR.n1480 2.04321
R2231 VDPWR.n1486 VDPWR.n1483 2.04321
R2232 VDPWR.n842 VDPWR.n781 2.04321
R2233 VDPWR.n941 VDPWR.n687 2.04321
R2234 VDPWR.n693 VDPWR.n690 2.04321
R2235 VDPWR.n934 VDPWR.n694 2.04321
R2236 VDPWR.n700 VDPWR.n697 2.04321
R2237 VDPWR.n927 VDPWR.n701 2.04321
R2238 VDPWR.n707 VDPWR.n704 2.04321
R2239 VDPWR.n920 VDPWR.n708 2.04321
R2240 VDPWR.n714 VDPWR.n711 2.04321
R2241 VDPWR.n913 VDPWR.n715 2.04321
R2242 VDPWR.n721 VDPWR.n718 2.04321
R2243 VDPWR.n906 VDPWR.n722 2.04321
R2244 VDPWR.n728 VDPWR.n725 2.04321
R2245 VDPWR.n899 VDPWR.n729 2.04321
R2246 VDPWR.n735 VDPWR.n732 2.04321
R2247 VDPWR.n892 VDPWR.n736 2.04321
R2248 VDPWR.n742 VDPWR.n739 2.04321
R2249 VDPWR.n885 VDPWR.n743 2.04321
R2250 VDPWR.n749 VDPWR.n746 2.04321
R2251 VDPWR.n878 VDPWR.n750 2.04321
R2252 VDPWR.n756 VDPWR.n753 2.04321
R2253 VDPWR.n871 VDPWR.n757 2.04321
R2254 VDPWR.n763 VDPWR.n760 2.04321
R2255 VDPWR.n864 VDPWR.n764 2.04321
R2256 VDPWR.n770 VDPWR.n767 2.04321
R2257 VDPWR.n857 VDPWR.n771 2.04321
R2258 VDPWR.n777 VDPWR.n774 2.04321
R2259 VDPWR.n850 VDPWR.n778 2.04321
R2260 VDPWR.n843 VDPWR.n841 2.04321
R2261 VDPWR.n477 VDPWR.n190 2.04321
R2262 VDPWR.n476 VDPWR.n189 2.04321
R2263 VDPWR.n183 VDPWR.n182 2.04321
R2264 VDPWR.n487 VDPWR.n181 2.04321
R2265 VDPWR.n451 VDPWR.n214 2.04321
R2266 VDPWR.n450 VDPWR.n213 2.04321
R2267 VDPWR.n207 VDPWR.n206 2.04321
R2268 VDPWR.n461 VDPWR.n205 2.04321
R2269 VDPWR.n425 VDPWR.n238 2.04321
R2270 VDPWR.n424 VDPWR.n237 2.04321
R2271 VDPWR.n231 VDPWR.n230 2.04321
R2272 VDPWR.n435 VDPWR.n229 2.04321
R2273 VDPWR.n399 VDPWR.n262 2.04321
R2274 VDPWR.n398 VDPWR.n261 2.04321
R2275 VDPWR.n255 VDPWR.n254 2.04321
R2276 VDPWR.n409 VDPWR.n253 2.04321
R2277 VDPWR.n373 VDPWR.n286 2.04321
R2278 VDPWR.n372 VDPWR.n285 2.04321
R2279 VDPWR.n279 VDPWR.n278 2.04321
R2280 VDPWR.n383 VDPWR.n277 2.04321
R2281 VDPWR.n339 VDPWR.n310 2.04321
R2282 VDPWR.n338 VDPWR.n309 2.04321
R2283 VDPWR.n303 VDPWR.n302 2.04321
R2284 VDPWR.n349 VDPWR.n301 2.04321
R2285 VDPWR.n108 VDPWR.n21 2.04321
R2286 VDPWR.n107 VDPWR.n20 2.04321
R2287 VDPWR.n14 VDPWR.n13 2.04321
R2288 VDPWR.n118 VDPWR.n12 2.04321
R2289 VDPWR.n74 VDPWR.n45 2.04321
R2290 VDPWR.n84 VDPWR.n36 2.04321
R2291 VDPWR.n38 VDPWR.n37 2.04321
R2292 VDPWR.n982 VDPWR.n981 1.97967
R2293 VDPWR.n1000 VDPWR.n999 1.97967
R2294 VDPWR.n1018 VDPWR.n1017 1.97967
R2295 VDPWR.n1036 VDPWR.n1035 1.97967
R2296 VDPWR.n1054 VDPWR.n1053 1.97967
R2297 VDPWR.n1072 VDPWR.n1071 1.97967
R2298 VDPWR.n1090 VDPWR.n1089 1.97967
R2299 VDPWR.n1108 VDPWR.n1107 1.97967
R2300 VDPWR VDPWR.n322 1.97234
R2301 VDPWR VDPWR.n57 1.97234
R2302 VDPWR.n491 VDPWR.n490 1.96588
R2303 VDPWR.n499 VDPWR.n175 1.96588
R2304 VDPWR.n502 VDPWR.n501 1.96588
R2305 VDPWR.n510 VDPWR.n169 1.96588
R2306 VDPWR.n130 VDPWR.n129 1.96588
R2307 VDPWR.n138 VDPWR.n6 1.96588
R2308 VDPWR.n141 VDPWR.n140 1.96588
R2309 VDPWR.n149 VDPWR.n0 1.96588
R2310 VDPWR.n466 VDPWR.n199 1.96583
R2311 VDPWR.n462 VDPWR.n202 1.96583
R2312 VDPWR.n195 VDPWR.n194 1.96583
R2313 VDPWR.n475 VDPWR.n191 1.96583
R2314 VDPWR.n440 VDPWR.n223 1.96583
R2315 VDPWR.n436 VDPWR.n226 1.96583
R2316 VDPWR.n219 VDPWR.n218 1.96583
R2317 VDPWR.n449 VDPWR.n215 1.96583
R2318 VDPWR.n414 VDPWR.n247 1.96583
R2319 VDPWR.n410 VDPWR.n250 1.96583
R2320 VDPWR.n243 VDPWR.n242 1.96583
R2321 VDPWR.n423 VDPWR.n239 1.96583
R2322 VDPWR.n388 VDPWR.n271 1.96583
R2323 VDPWR.n384 VDPWR.n274 1.96583
R2324 VDPWR.n267 VDPWR.n266 1.96583
R2325 VDPWR.n397 VDPWR.n263 1.96583
R2326 VDPWR.n362 VDPWR.n295 1.96583
R2327 VDPWR.n358 VDPWR.n298 1.96583
R2328 VDPWR.n291 VDPWR.n290 1.96583
R2329 VDPWR.n371 VDPWR.n287 1.96583
R2330 VDPWR.n328 VDPWR.n319 1.96583
R2331 VDPWR.n315 VDPWR.n314 1.96583
R2332 VDPWR.n337 VDPWR.n311 1.96583
R2333 VDPWR.n97 VDPWR.n30 1.96583
R2334 VDPWR.n93 VDPWR.n33 1.96583
R2335 VDPWR.n26 VDPWR.n25 1.96583
R2336 VDPWR.n106 VDPWR.n22 1.96583
R2337 VDPWR.n63 VDPWR.n54 1.96583
R2338 VDPWR.n50 VDPWR.n49 1.96583
R2339 VDPWR.n72 VDPWR.n46 1.96583
R2340 VDPWR.n1180 VDPWR.n1159 1.9397
R2341 VDPWR.n1184 VDPWR.n1183 1.9397
R2342 VDPWR.n1196 VDPWR.n1154 1.9397
R2343 VDPWR.n1200 VDPWR.n1199 1.9397
R2344 VDPWR.n1212 VDPWR.n1149 1.9397
R2345 VDPWR.n1216 VDPWR.n1215 1.9397
R2346 VDPWR.n1228 VDPWR.n1144 1.9397
R2347 VDPWR.n1232 VDPWR.n1231 1.9397
R2348 VDPWR.n1244 VDPWR.n1139 1.9397
R2349 VDPWR.n1248 VDPWR.n1247 1.9397
R2350 VDPWR.n1260 VDPWR.n1134 1.9397
R2351 VDPWR.n1264 VDPWR.n1263 1.9397
R2352 VDPWR.n1276 VDPWR.n1129 1.9397
R2353 VDPWR.n1280 VDPWR.n1279 1.9397
R2354 VDPWR.n1292 VDPWR.n1124 1.9397
R2355 VDPWR.n1296 VDPWR.n1295 1.9397
R2356 VDPWR.n1308 VDPWR.n1119 1.9397
R2357 VDPWR.n1385 VDPWR.n1359 1.9397
R2358 VDPWR.n1386 VDPWR.n1355 1.9397
R2359 VDPWR.n1395 VDPWR.n1354 1.9397
R2360 VDPWR.n1353 VDPWR.n1348 1.9397
R2361 VDPWR.n1413 VDPWR.n1343 1.9397
R2362 VDPWR.n1414 VDPWR.n1339 1.9397
R2363 VDPWR.n1423 VDPWR.n1338 1.9397
R2364 VDPWR.n1337 VDPWR.n1332 1.9397
R2365 VDPWR.n1441 VDPWR.n1327 1.9397
R2366 VDPWR.n1442 VDPWR.n1323 1.9397
R2367 VDPWR.n1451 VDPWR.n1322 1.9397
R2368 VDPWR.n1321 VDPWR.n1316 1.9397
R2369 VDPWR.n1465 VDPWR.n1311 1.9397
R2370 VDPWR.n165 VDPWR.n163 1.8605
R2371 VDPWR.n179 VDPWR.n176 1.54255
R2372 VDPWR.n173 VDPWR.n170 1.54255
R2373 VDPWR.n10 VDPWR.n7 1.54255
R2374 VDPWR.n4 VDPWR.n1 1.54255
R2375 VDPWR.n1183 VDPWR.n1180 1.52654
R2376 VDPWR.n1199 VDPWR.n1196 1.52654
R2377 VDPWR.n1215 VDPWR.n1212 1.52654
R2378 VDPWR.n1231 VDPWR.n1228 1.52654
R2379 VDPWR.n1247 VDPWR.n1244 1.52654
R2380 VDPWR.n1263 VDPWR.n1260 1.52654
R2381 VDPWR.n1279 VDPWR.n1276 1.52654
R2382 VDPWR.n1295 VDPWR.n1292 1.52654
R2383 VDPWR.n681 VDPWR.n677 1.51949
R2384 VDPWR.n664 VDPWR.n660 1.51949
R2385 VDPWR.n647 VDPWR.n643 1.51949
R2386 VDPWR.n630 VDPWR.n626 1.51949
R2387 VDPWR.n613 VDPWR.n609 1.51949
R2388 VDPWR.n596 VDPWR.n592 1.51949
R2389 VDPWR.n579 VDPWR.n575 1.51949
R2390 VDPWR.n562 VDPWR.n558 1.51949
R2391 VDPWR.n1545 VDPWR.n1544 1.45922
R2392 VDPWR.n1309 VDPWR.n1118 1.39972
R2393 VDPWR.n129 VDPWR 1.37724
R2394 VDPWR.n335 VDPWR.n334 1.32907
R2395 VDPWR.n327 VDPWR.n326 1.32907
R2396 VDPWR.n369 VDPWR.n368 1.32907
R2397 VDPWR.n361 VDPWR.n360 1.32907
R2398 VDPWR.n395 VDPWR.n394 1.32907
R2399 VDPWR.n387 VDPWR.n386 1.32907
R2400 VDPWR.n421 VDPWR.n420 1.32907
R2401 VDPWR.n413 VDPWR.n412 1.32907
R2402 VDPWR.n447 VDPWR.n446 1.32907
R2403 VDPWR.n439 VDPWR.n438 1.32907
R2404 VDPWR.n473 VDPWR.n472 1.32907
R2405 VDPWR.n465 VDPWR.n464 1.32907
R2406 VDPWR.n70 VDPWR.n69 1.32907
R2407 VDPWR.n62 VDPWR.n61 1.32907
R2408 VDPWR.n104 VDPWR.n103 1.32907
R2409 VDPWR.n96 VDPWR.n95 1.32907
R2410 VDPWR.n354 VDPWR 1.24128
R2411 VDPWR.n123 VDPWR 1.24128
R2412 VDPWR.n89 VDPWR 1.24128
R2413 VDPWR.n490 VDPWR 1.23314
R2414 VDPWR.n463 VDPWR.n204 1.21789
R2415 VDPWR.n474 VDPWR.n193 1.21789
R2416 VDPWR.n437 VDPWR.n228 1.21789
R2417 VDPWR.n448 VDPWR.n217 1.21789
R2418 VDPWR.n411 VDPWR.n252 1.21789
R2419 VDPWR.n422 VDPWR.n241 1.21789
R2420 VDPWR.n385 VDPWR.n276 1.21789
R2421 VDPWR.n396 VDPWR.n265 1.21789
R2422 VDPWR.n359 VDPWR.n300 1.21789
R2423 VDPWR.n370 VDPWR.n289 1.21789
R2424 VDPWR.n325 VDPWR.n324 1.21789
R2425 VDPWR.n336 VDPWR.n313 1.21789
R2426 VDPWR.n94 VDPWR.n35 1.21789
R2427 VDPWR.n105 VDPWR.n24 1.21789
R2428 VDPWR.n60 VDPWR.n59 1.21789
R2429 VDPWR.n71 VDPWR.n48 1.21789
R2430 VDPWR.n1192 VDPWR.n1191 1.21332
R2431 VDPWR.n1208 VDPWR.n1207 1.21332
R2432 VDPWR.n1224 VDPWR.n1223 1.21332
R2433 VDPWR.n1240 VDPWR.n1239 1.21332
R2434 VDPWR.n1256 VDPWR.n1255 1.21332
R2435 VDPWR.n1272 VDPWR.n1271 1.21332
R2436 VDPWR.n1288 VDPWR.n1287 1.21332
R2437 VDPWR.n1304 VDPWR.n1303 1.21332
R2438 VDPWR.n1394 VDPWR.n1356 1.21332
R2439 VDPWR.n1409 VDPWR.n1408 1.21332
R2440 VDPWR.n1422 VDPWR.n1340 1.21332
R2441 VDPWR.n1437 VDPWR.n1436 1.21332
R2442 VDPWR.n1450 VDPWR.n1324 1.21332
R2443 VDPWR.n1461 VDPWR.n1460 1.21332
R2444 VDPWR.n352 VDPWR.n351 1.09595
R2445 VDPWR.n121 VDPWR.n120 1.09595
R2446 VDPWR.n87 VDPWR.n86 1.09595
R2447 VDPWR.n568 VDPWR 1.04243
R2448 VDPWR.n585 VDPWR 1.04243
R2449 VDPWR.n602 VDPWR 1.04243
R2450 VDPWR.n619 VDPWR 1.04243
R2451 VDPWR.n636 VDPWR 1.04243
R2452 VDPWR.n653 VDPWR 1.04243
R2453 VDPWR.n670 VDPWR 1.04243
R2454 VDPWR.n1117 VDPWR.n941 0.948417
R2455 VDPWR.n548 VDPWR.n547 0.832022
R2456 VDPWR.n543 VDPWR.n542 0.832022
R2457 VDPWR.n538 VDPWR.n537 0.832022
R2458 VDPWR.n533 VDPWR.n532 0.832022
R2459 VDPWR.n528 VDPWR.n527 0.832022
R2460 VDPWR.n523 VDPWR.n522 0.832022
R2461 VDPWR.n518 VDPWR.n517 0.832022
R2462 VDPWR.n513 VDPWR.n512 0.832022
R2463 VDPWR VDPWR.n1308 0.813
R2464 VDPWR.n356 VDPWR.n355 0.8005
R2465 VDPWR.n91 VDPWR.n90 0.795143
R2466 VDPWR.n125 VDPWR.n124 0.777286
R2467 VDPWR.n127 VDPWR 0.7505
R2468 VDPWR.n1543 VDPWR.n1542 0.68153
R2469 VDPWR.n993 VDPWR 0.669618
R2470 VDPWR.n1011 VDPWR 0.669618
R2471 VDPWR.n1029 VDPWR 0.669618
R2472 VDPWR.n1047 VDPWR 0.669618
R2473 VDPWR.n1065 VDPWR 0.669618
R2474 VDPWR.n1083 VDPWR 0.669618
R2475 VDPWR.n1101 VDPWR 0.669618
R2476 VDPWR.n161 VDPWR.n150 0.6555
R2477 VDPWR.n552 VDPWR.n550 0.629553
R2478 VDPWR.n1305 VDPWR.n1304 0.6205
R2479 VDPWR.n1289 VDPWR.n1288 0.6205
R2480 VDPWR.n1273 VDPWR.n1272 0.6205
R2481 VDPWR.n1257 VDPWR.n1256 0.6205
R2482 VDPWR.n1241 VDPWR.n1240 0.6205
R2483 VDPWR.n1225 VDPWR.n1224 0.6205
R2484 VDPWR.n1209 VDPWR.n1208 0.6205
R2485 VDPWR.n1193 VDPWR.n1192 0.6205
R2486 VDPWR.n1177 VDPWR.n1176 0.6205
R2487 VDPWR.n1462 VDPWR.n1461 0.6205
R2488 VDPWR.n1450 VDPWR.n1449 0.6205
R2489 VDPWR.n1438 VDPWR.n1437 0.6205
R2490 VDPWR.n1422 VDPWR.n1421 0.6205
R2491 VDPWR.n1410 VDPWR.n1409 0.6205
R2492 VDPWR.n1394 VDPWR.n1393 0.6205
R2493 VDPWR.n1382 VDPWR.n1381 0.6205
R2494 VDPWR.n550 VDPWR.n549 0.61463
R2495 VDPWR.n545 VDPWR.n544 0.61463
R2496 VDPWR.n540 VDPWR.n539 0.61463
R2497 VDPWR.n535 VDPWR.n534 0.61463
R2498 VDPWR.n530 VDPWR.n529 0.61463
R2499 VDPWR.n525 VDPWR.n524 0.61463
R2500 VDPWR.n520 VDPWR.n519 0.61463
R2501 VDPWR.n515 VDPWR.n514 0.61463
R2502 VDPWR.n1551 VDPWR.n161 0.60099
R2503 VDPWR.n1112 VDPWR.n1111 0.58175
R2504 VDPWR.n1094 VDPWR.n1093 0.58175
R2505 VDPWR.n1076 VDPWR.n1075 0.58175
R2506 VDPWR.n1058 VDPWR.n1057 0.58175
R2507 VDPWR.n1040 VDPWR.n1039 0.58175
R2508 VDPWR.n1022 VDPWR.n1021 0.58175
R2509 VDPWR.n1004 VDPWR.n1003 0.58175
R2510 VDPWR.n986 VDPWR.n985 0.58175
R2511 VDPWR VDPWR.n383 0.568208
R2512 VDPWR VDPWR.n409 0.568208
R2513 VDPWR VDPWR.n435 0.568208
R2514 VDPWR VDPWR.n461 0.568208
R2515 VDPWR.n1176 VDPWR.n1164 0.533833
R2516 VDPWR.n1381 VDPWR.n1364 0.533833
R2517 VDPWR.n150 VDPWR 0.472722
R2518 VDPWR.n501 VDPWR 0.453625
R2519 VDPWR.n140 VDPWR 0.453625
R2520 VDPWR.n338 VDPWR 0.432792
R2521 VDPWR.n372 VDPWR 0.432792
R2522 VDPWR.n398 VDPWR 0.432792
R2523 VDPWR.n424 VDPWR 0.432792
R2524 VDPWR.n450 VDPWR 0.432792
R2525 VDPWR.n476 VDPWR 0.432792
R2526 VDPWR.n107 VDPWR 0.432792
R2527 VDPWR.n319 VDPWR.n314 0.430188
R2528 VDPWR.n295 VDPWR.n290 0.430188
R2529 VDPWR.n271 VDPWR.n266 0.430188
R2530 VDPWR.n247 VDPWR.n242 0.430188
R2531 VDPWR.n223 VDPWR.n218 0.430188
R2532 VDPWR.n199 VDPWR.n194 0.430188
R2533 VDPWR.n54 VDPWR.n49 0.430188
R2534 VDPWR.n30 VDPWR.n25 0.430188
R2535 VDPWR.n508 VDPWR.n507 0.423227
R2536 VDPWR.n497 VDPWR.n496 0.423227
R2537 VDPWR.n147 VDPWR.n146 0.423227
R2538 VDPWR.n136 VDPWR.n135 0.423227
R2539 VDPWR.n354 VDPWR 0.402286
R2540 VDPWR.n123 VDPWR 0.402286
R2541 VDPWR.n89 VDPWR 0.402286
R2542 VDPWR.n73 VDPWR 0.401542
R2543 VDPWR.n1543 VDPWR 0.392832
R2544 VDPWR VDPWR.n357 0.389823
R2545 VDPWR VDPWR.n92 0.385917
R2546 VDPWR VDPWR.n567 0.3755
R2547 VDPWR VDPWR.n584 0.3755
R2548 VDPWR VDPWR.n601 0.3755
R2549 VDPWR VDPWR.n618 0.3755
R2550 VDPWR VDPWR.n635 0.3755
R2551 VDPWR VDPWR.n652 0.3755
R2552 VDPWR VDPWR.n669 0.3755
R2553 VDPWR VDPWR.n686 0.3755
R2554 VDPWR.n326 VDPWR.n319 0.359875
R2555 VDPWR.n335 VDPWR.n314 0.359875
R2556 VDPWR.n360 VDPWR.n295 0.359875
R2557 VDPWR.n369 VDPWR.n290 0.359875
R2558 VDPWR.n386 VDPWR.n271 0.359875
R2559 VDPWR.n395 VDPWR.n266 0.359875
R2560 VDPWR.n412 VDPWR.n247 0.359875
R2561 VDPWR.n421 VDPWR.n242 0.359875
R2562 VDPWR.n438 VDPWR.n223 0.359875
R2563 VDPWR.n447 VDPWR.n218 0.359875
R2564 VDPWR.n464 VDPWR.n199 0.359875
R2565 VDPWR.n473 VDPWR.n194 0.359875
R2566 VDPWR.n61 VDPWR.n54 0.359875
R2567 VDPWR.n70 VDPWR.n49 0.359875
R2568 VDPWR.n95 VDPWR.n30 0.359875
R2569 VDPWR.n104 VDPWR.n25 0.359875
R2570 VDPWR.n569 VDPWR.n568 0.358192
R2571 VDPWR.n586 VDPWR.n585 0.358192
R2572 VDPWR.n603 VDPWR.n602 0.358192
R2573 VDPWR.n620 VDPWR.n619 0.358192
R2574 VDPWR.n637 VDPWR.n636 0.358192
R2575 VDPWR.n654 VDPWR.n653 0.358192
R2576 VDPWR.n671 VDPWR.n670 0.358192
R2577 VDPWR.n488 VDPWR.n487 0.357271
R2578 VDPWR.n549 VDPWR.n548 0.353761
R2579 VDPWR.n544 VDPWR.n543 0.353761
R2580 VDPWR.n539 VDPWR.n538 0.353761
R2581 VDPWR.n534 VDPWR.n533 0.353761
R2582 VDPWR.n529 VDPWR.n528 0.353761
R2583 VDPWR.n524 VDPWR.n523 0.353761
R2584 VDPWR.n519 VDPWR.n518 0.353761
R2585 VDPWR.n514 VDPWR.n513 0.353761
R2586 VDPWR.n1118 VDPWR 0.350184
R2587 VDPWR.n488 VDPWR 0.333833
R2588 VDPWR.n975 VDPWR.n973 0.324029
R2589 VDPWR.n989 VDPWR.n988 0.324029
R2590 VDPWR.n992 VDPWR.n969 0.324029
R2591 VDPWR.n1007 VDPWR.n1006 0.324029
R2592 VDPWR.n1010 VDPWR.n965 0.324029
R2593 VDPWR.n1025 VDPWR.n1024 0.324029
R2594 VDPWR.n1028 VDPWR.n961 0.324029
R2595 VDPWR.n1043 VDPWR.n1042 0.324029
R2596 VDPWR.n1046 VDPWR.n957 0.324029
R2597 VDPWR.n1061 VDPWR.n1060 0.324029
R2598 VDPWR.n1064 VDPWR.n953 0.324029
R2599 VDPWR.n1079 VDPWR.n1078 0.324029
R2600 VDPWR.n1082 VDPWR.n949 0.324029
R2601 VDPWR.n1097 VDPWR.n1096 0.324029
R2602 VDPWR.n1100 VDPWR.n945 0.324029
R2603 VDPWR.n1115 VDPWR.n1114 0.324029
R2604 VDPWR.n1118 VDPWR.n1117 0.274719
R2605 VDPWR.n568 VDPWR.n545 0.271861
R2606 VDPWR.n585 VDPWR.n540 0.271861
R2607 VDPWR.n602 VDPWR.n535 0.271861
R2608 VDPWR.n619 VDPWR.n530 0.271861
R2609 VDPWR.n636 VDPWR.n525 0.271861
R2610 VDPWR.n653 VDPWR.n520 0.271861
R2611 VDPWR.n670 VDPWR.n515 0.271861
R2612 VDPWR.n1177 VDPWR.n1163 0.253104
R2613 VDPWR.n1193 VDPWR.n1158 0.253104
R2614 VDPWR.n1209 VDPWR.n1153 0.253104
R2615 VDPWR.n1225 VDPWR.n1148 0.253104
R2616 VDPWR.n1241 VDPWR.n1143 0.253104
R2617 VDPWR.n1257 VDPWR.n1138 0.253104
R2618 VDPWR.n1273 VDPWR.n1133 0.253104
R2619 VDPWR.n1289 VDPWR.n1128 0.253104
R2620 VDPWR.n1305 VDPWR.n1123 0.253104
R2621 VDPWR.n1382 VDPWR.n1363 0.253104
R2622 VDPWR.n1393 VDPWR.n1388 0.253104
R2623 VDPWR.n1410 VDPWR.n1347 0.253104
R2624 VDPWR.n1421 VDPWR.n1416 0.253104
R2625 VDPWR.n1438 VDPWR.n1331 0.253104
R2626 VDPWR.n1449 VDPWR.n1444 0.253104
R2627 VDPWR.n1462 VDPWR.n1315 0.253104
R2628 VDPWR.n985 VDPWR.n984 0.25148
R2629 VDPWR.n1003 VDPWR.n1002 0.25148
R2630 VDPWR.n1021 VDPWR.n1020 0.25148
R2631 VDPWR.n1039 VDPWR.n1038 0.25148
R2632 VDPWR.n1057 VDPWR.n1056 0.25148
R2633 VDPWR.n1075 VDPWR.n1074 0.25148
R2634 VDPWR.n1093 VDPWR.n1092 0.25148
R2635 VDPWR.n1111 VDPWR.n1110 0.25148
R2636 VDPWR.n1180 VDPWR.n1179 0.246594
R2637 VDPWR.n1183 VDPWR.n1182 0.246594
R2638 VDPWR.n1196 VDPWR.n1195 0.246594
R2639 VDPWR.n1199 VDPWR.n1198 0.246594
R2640 VDPWR.n1212 VDPWR.n1211 0.246594
R2641 VDPWR.n1215 VDPWR.n1214 0.246594
R2642 VDPWR.n1228 VDPWR.n1227 0.246594
R2643 VDPWR.n1231 VDPWR.n1230 0.246594
R2644 VDPWR.n1244 VDPWR.n1243 0.246594
R2645 VDPWR.n1247 VDPWR.n1246 0.246594
R2646 VDPWR.n1260 VDPWR.n1259 0.246594
R2647 VDPWR.n1263 VDPWR.n1262 0.246594
R2648 VDPWR.n1276 VDPWR.n1275 0.246594
R2649 VDPWR.n1279 VDPWR.n1278 0.246594
R2650 VDPWR.n1292 VDPWR.n1291 0.246594
R2651 VDPWR.n1295 VDPWR.n1294 0.246594
R2652 VDPWR.n1308 VDPWR.n1307 0.246594
R2653 VDPWR.n1385 VDPWR.n1384 0.246594
R2654 VDPWR.n1387 VDPWR.n1386 0.246594
R2655 VDPWR.n1391 VDPWR.n1354 0.246594
R2656 VDPWR.n1353 VDPWR.n1352 0.246594
R2657 VDPWR.n1413 VDPWR.n1412 0.246594
R2658 VDPWR.n1415 VDPWR.n1414 0.246594
R2659 VDPWR.n1419 VDPWR.n1338 0.246594
R2660 VDPWR.n1337 VDPWR.n1336 0.246594
R2661 VDPWR.n1441 VDPWR.n1440 0.246594
R2662 VDPWR.n1443 VDPWR.n1442 0.246594
R2663 VDPWR.n1447 VDPWR.n1322 0.246594
R2664 VDPWR.n1321 VDPWR.n1320 0.246594
R2665 VDPWR.n1465 VDPWR.n1464 0.246594
R2666 VDPWR.n1178 VDPWR.n1177 0.242688
R2667 VDPWR.n1194 VDPWR.n1193 0.242688
R2668 VDPWR.n1210 VDPWR.n1209 0.242688
R2669 VDPWR.n1226 VDPWR.n1225 0.242688
R2670 VDPWR.n1242 VDPWR.n1241 0.242688
R2671 VDPWR.n1258 VDPWR.n1257 0.242688
R2672 VDPWR.n1274 VDPWR.n1273 0.242688
R2673 VDPWR.n1290 VDPWR.n1289 0.242688
R2674 VDPWR.n1306 VDPWR.n1305 0.242688
R2675 VDPWR.n1383 VDPWR.n1382 0.242688
R2676 VDPWR.n1393 VDPWR.n1392 0.242688
R2677 VDPWR.n1411 VDPWR.n1410 0.242688
R2678 VDPWR.n1421 VDPWR.n1420 0.242688
R2679 VDPWR.n1439 VDPWR.n1438 0.242688
R2680 VDPWR.n1449 VDPWR.n1448 0.242688
R2681 VDPWR.n1463 VDPWR.n1462 0.242688
R2682 VDPWR.n511 VDPWR 0.241819
R2683 VDPWR.n1541 VDPWR 0.240083
R2684 VDPWR.n993 VDPWR.n992 0.239471
R2685 VDPWR.n1011 VDPWR.n1010 0.239471
R2686 VDPWR.n1029 VDPWR.n1028 0.239471
R2687 VDPWR.n1047 VDPWR.n1046 0.239471
R2688 VDPWR.n1065 VDPWR.n1064 0.239471
R2689 VDPWR.n1083 VDPWR.n1082 0.239471
R2690 VDPWR.n1101 VDPWR.n1100 0.239471
R2691 VDPWR.n990 VDPWR.n989 0.232118
R2692 VDPWR.n1008 VDPWR.n1007 0.232118
R2693 VDPWR.n1026 VDPWR.n1025 0.232118
R2694 VDPWR.n1044 VDPWR.n1043 0.232118
R2695 VDPWR.n1062 VDPWR.n1061 0.232118
R2696 VDPWR.n1080 VDPWR.n1079 0.232118
R2697 VDPWR.n1098 VDPWR.n1097 0.232118
R2698 VDPWR.n1116 VDPWR.n1115 0.232118
R2699 VDPWR.n1168 VDPWR.n1163 0.229667
R2700 VDPWR.n1179 VDPWR.n1178 0.229667
R2701 VDPWR.n1182 VDPWR.n1158 0.229667
R2702 VDPWR.n1195 VDPWR.n1194 0.229667
R2703 VDPWR.n1198 VDPWR.n1153 0.229667
R2704 VDPWR.n1211 VDPWR.n1210 0.229667
R2705 VDPWR.n1214 VDPWR.n1148 0.229667
R2706 VDPWR.n1227 VDPWR.n1226 0.229667
R2707 VDPWR.n1230 VDPWR.n1143 0.229667
R2708 VDPWR.n1243 VDPWR.n1242 0.229667
R2709 VDPWR.n1246 VDPWR.n1138 0.229667
R2710 VDPWR.n1259 VDPWR.n1258 0.229667
R2711 VDPWR.n1262 VDPWR.n1133 0.229667
R2712 VDPWR.n1275 VDPWR.n1274 0.229667
R2713 VDPWR.n1278 VDPWR.n1128 0.229667
R2714 VDPWR.n1291 VDPWR.n1290 0.229667
R2715 VDPWR.n1294 VDPWR.n1123 0.229667
R2716 VDPWR.n1307 VDPWR.n1306 0.229667
R2717 VDPWR.n1384 VDPWR.n1383 0.229667
R2718 VDPWR.n1388 VDPWR.n1387 0.229667
R2719 VDPWR.n1392 VDPWR.n1391 0.229667
R2720 VDPWR.n1352 VDPWR.n1347 0.229667
R2721 VDPWR.n1412 VDPWR.n1411 0.229667
R2722 VDPWR.n1416 VDPWR.n1415 0.229667
R2723 VDPWR.n1420 VDPWR.n1419 0.229667
R2724 VDPWR.n1336 VDPWR.n1331 0.229667
R2725 VDPWR.n1440 VDPWR.n1439 0.229667
R2726 VDPWR.n1444 VDPWR.n1443 0.229667
R2727 VDPWR.n1448 VDPWR.n1447 0.229667
R2728 VDPWR.n1320 VDPWR.n1315 0.229667
R2729 VDPWR.n1464 VDPWR.n1463 0.229667
R2730 VDPWR.n326 VDPWR.n325 0.229667
R2731 VDPWR.n336 VDPWR.n335 0.229667
R2732 VDPWR.n360 VDPWR.n359 0.229667
R2733 VDPWR.n370 VDPWR.n369 0.229667
R2734 VDPWR.n386 VDPWR.n385 0.229667
R2735 VDPWR.n396 VDPWR.n395 0.229667
R2736 VDPWR.n412 VDPWR.n411 0.229667
R2737 VDPWR.n422 VDPWR.n421 0.229667
R2738 VDPWR.n438 VDPWR.n437 0.229667
R2739 VDPWR.n448 VDPWR.n447 0.229667
R2740 VDPWR.n464 VDPWR.n463 0.229667
R2741 VDPWR.n474 VDPWR.n473 0.229667
R2742 VDPWR.n61 VDPWR.n60 0.229667
R2743 VDPWR.n71 VDPWR.n70 0.229667
R2744 VDPWR.n95 VDPWR.n94 0.229667
R2745 VDPWR.n105 VDPWR.n104 0.229667
R2746 VDPWR.n161 VDPWR.n160 0.223
R2747 VDPWR.n1386 VDPWR.n1385 0.221854
R2748 VDPWR.n1354 VDPWR.n1353 0.221854
R2749 VDPWR.n1414 VDPWR.n1413 0.221854
R2750 VDPWR.n1338 VDPWR.n1337 0.221854
R2751 VDPWR.n1442 VDPWR.n1441 0.221854
R2752 VDPWR.n1322 VDPWR.n1321 0.221854
R2753 VDPWR.n1509 VDPWR 0.2005
R2754 VDPWR.n1368 VDPWR.n1363 0.199719
R2755 VDPWR.n126 VDPWR.n118 0.195812
R2756 VDPWR.n941 VDPWR.n940 0.189302
R2757 VDPWR.n936 VDPWR.n693 0.189302
R2758 VDPWR.n934 VDPWR.n933 0.189302
R2759 VDPWR.n929 VDPWR.n700 0.189302
R2760 VDPWR.n927 VDPWR.n926 0.189302
R2761 VDPWR.n922 VDPWR.n707 0.189302
R2762 VDPWR.n920 VDPWR.n919 0.189302
R2763 VDPWR.n915 VDPWR.n714 0.189302
R2764 VDPWR.n913 VDPWR.n912 0.189302
R2765 VDPWR.n908 VDPWR.n721 0.189302
R2766 VDPWR.n906 VDPWR.n905 0.189302
R2767 VDPWR.n901 VDPWR.n728 0.189302
R2768 VDPWR.n899 VDPWR.n898 0.189302
R2769 VDPWR.n894 VDPWR.n735 0.189302
R2770 VDPWR.n892 VDPWR.n891 0.189302
R2771 VDPWR.n887 VDPWR.n742 0.189302
R2772 VDPWR.n885 VDPWR.n884 0.189302
R2773 VDPWR.n880 VDPWR.n749 0.189302
R2774 VDPWR.n878 VDPWR.n877 0.189302
R2775 VDPWR.n873 VDPWR.n756 0.189302
R2776 VDPWR.n871 VDPWR.n870 0.189302
R2777 VDPWR.n866 VDPWR.n763 0.189302
R2778 VDPWR.n864 VDPWR.n863 0.189302
R2779 VDPWR.n859 VDPWR.n770 0.189302
R2780 VDPWR.n857 VDPWR.n856 0.189302
R2781 VDPWR.n852 VDPWR.n777 0.189302
R2782 VDPWR.n850 VDPWR.n849 0.189302
R2783 VDPWR.n845 VDPWR.n842 0.189302
R2784 VDPWR.n1540 VDPWR.n1539 0.189302
R2785 VDPWR.n1535 VDPWR.n1472 0.189302
R2786 VDPWR.n1533 VDPWR.n1532 0.189302
R2787 VDPWR.n1528 VDPWR.n1479 0.189302
R2788 VDPWR.n1526 VDPWR.n1525 0.189302
R2789 VDPWR.n1521 VDPWR.n1486 0.189302
R2790 VDPWR.n341 VDPWR.n338 0.189302
R2791 VDPWR.n347 VDPWR.n302 0.189302
R2792 VDPWR.n375 VDPWR.n372 0.189302
R2793 VDPWR.n381 VDPWR.n278 0.189302
R2794 VDPWR.n401 VDPWR.n398 0.189302
R2795 VDPWR.n407 VDPWR.n254 0.189302
R2796 VDPWR.n427 VDPWR.n424 0.189302
R2797 VDPWR.n433 VDPWR.n230 0.189302
R2798 VDPWR.n453 VDPWR.n450 0.189302
R2799 VDPWR.n459 VDPWR.n206 0.189302
R2800 VDPWR.n479 VDPWR.n476 0.189302
R2801 VDPWR.n485 VDPWR.n182 0.189302
R2802 VDPWR.n82 VDPWR.n37 0.189302
R2803 VDPWR.n110 VDPWR.n107 0.189302
R2804 VDPWR.n116 VDPWR.n13 0.189302
R2805 VDPWR.n1369 VDPWR.n1368 0.185396
R2806 VDPWR VDPWR.n499 0.182792
R2807 VDPWR VDPWR.n510 0.182792
R2808 VDPWR.n92 VDPWR.n84 0.182792
R2809 VDPWR VDPWR.n138 0.182792
R2810 VDPWR VDPWR.n149 0.182792
R2811 VDPWR.n357 VDPWR.n349 0.178885
R2812 VDPWR.n1369 VDPWR.n1310 0.174979
R2813 VDPWR.n127 VDPWR.n126 0.174979
R2814 VDPWR.n490 VDPWR.n489 0.166299
R2815 VDPWR.n501 VDPWR.n500 0.166299
R2816 VDPWR.n129 VDPWR.n128 0.166299
R2817 VDPWR.n140 VDPWR.n139 0.166299
R2818 VDPWR.n1310 VDPWR 0.164562
R2819 VDPWR.n1519 VDPWR.n1487 0.158052
R2820 VDPWR.n1511 VDPWR.n1504 0.158052
R2821 VDPWR.n76 VDPWR.n73 0.158052
R2822 VDPWR VDPWR.n1465 0.151542
R2823 VDPWR.n339 VDPWR.n302 0.141125
R2824 VDPWR.n373 VDPWR.n278 0.141125
R2825 VDPWR.n399 VDPWR.n254 0.141125
R2826 VDPWR.n425 VDPWR.n230 0.141125
R2827 VDPWR.n451 VDPWR.n206 0.141125
R2828 VDPWR.n477 VDPWR.n182 0.141125
R2829 VDPWR.n74 VDPWR.n37 0.141125
R2830 VDPWR.n108 VDPWR.n13 0.141125
R2831 VDPWR VDPWR.n1551 0.133312
R2832 VDPWR.n693 VDPWR.n688 0.13201
R2833 VDPWR.n935 VDPWR.n934 0.13201
R2834 VDPWR.n700 VDPWR.n695 0.13201
R2835 VDPWR.n928 VDPWR.n927 0.13201
R2836 VDPWR.n707 VDPWR.n702 0.13201
R2837 VDPWR.n921 VDPWR.n920 0.13201
R2838 VDPWR.n714 VDPWR.n709 0.13201
R2839 VDPWR.n914 VDPWR.n913 0.13201
R2840 VDPWR.n721 VDPWR.n716 0.13201
R2841 VDPWR.n907 VDPWR.n906 0.13201
R2842 VDPWR.n728 VDPWR.n723 0.13201
R2843 VDPWR.n900 VDPWR.n899 0.13201
R2844 VDPWR.n735 VDPWR.n730 0.13201
R2845 VDPWR.n893 VDPWR.n892 0.13201
R2846 VDPWR.n742 VDPWR.n737 0.13201
R2847 VDPWR.n886 VDPWR.n885 0.13201
R2848 VDPWR.n749 VDPWR.n744 0.13201
R2849 VDPWR.n879 VDPWR.n878 0.13201
R2850 VDPWR.n756 VDPWR.n751 0.13201
R2851 VDPWR.n872 VDPWR.n871 0.13201
R2852 VDPWR.n763 VDPWR.n758 0.13201
R2853 VDPWR.n865 VDPWR.n864 0.13201
R2854 VDPWR.n770 VDPWR.n765 0.13201
R2855 VDPWR.n858 VDPWR.n857 0.13201
R2856 VDPWR.n777 VDPWR.n772 0.13201
R2857 VDPWR.n851 VDPWR.n850 0.13201
R2858 VDPWR.n842 VDPWR.n779 0.13201
R2859 VDPWR.n844 VDPWR.n843 0.13201
R2860 VDPWR.n1472 VDPWR.n1467 0.13201
R2861 VDPWR.n1534 VDPWR.n1533 0.13201
R2862 VDPWR.n1479 VDPWR.n1474 0.13201
R2863 VDPWR.n1527 VDPWR.n1526 0.13201
R2864 VDPWR.n1486 VDPWR.n1481 0.13201
R2865 VDPWR.n340 VDPWR.n339 0.13201
R2866 VDPWR.n349 VDPWR.n348 0.13201
R2867 VDPWR.n374 VDPWR.n373 0.13201
R2868 VDPWR.n383 VDPWR.n382 0.13201
R2869 VDPWR.n400 VDPWR.n399 0.13201
R2870 VDPWR.n409 VDPWR.n408 0.13201
R2871 VDPWR.n426 VDPWR.n425 0.13201
R2872 VDPWR.n435 VDPWR.n434 0.13201
R2873 VDPWR.n452 VDPWR.n451 0.13201
R2874 VDPWR.n461 VDPWR.n460 0.13201
R2875 VDPWR.n478 VDPWR.n477 0.13201
R2876 VDPWR.n487 VDPWR.n486 0.13201
R2877 VDPWR.n75 VDPWR.n74 0.13201
R2878 VDPWR.n84 VDPWR.n83 0.13201
R2879 VDPWR.n109 VDPWR.n108 0.13201
R2880 VDPWR.n118 VDPWR.n117 0.13201
R2881 VDPWR.n337 VDPWR.n336 0.130708
R2882 VDPWR.n371 VDPWR.n370 0.130708
R2883 VDPWR.n397 VDPWR.n396 0.130708
R2884 VDPWR.n423 VDPWR.n422 0.130708
R2885 VDPWR.n449 VDPWR.n448 0.130708
R2886 VDPWR.n475 VDPWR.n474 0.130708
R2887 VDPWR.n72 VDPWR.n71 0.130708
R2888 VDPWR.n106 VDPWR.n105 0.130708
R2889 VDPWR.n498 VDPWR.n497 0.127236
R2890 VDPWR.n509 VDPWR.n508 0.127236
R2891 VDPWR.n137 VDPWR.n136 0.127236
R2892 VDPWR.n148 VDPWR.n147 0.127236
R2893 VDPWR.n1509 VDPWR 0.1255
R2894 VDPWR.n988 VDPWR.n987 0.124275
R2895 VDPWR.n1006 VDPWR.n1005 0.124275
R2896 VDPWR.n1024 VDPWR.n1023 0.124275
R2897 VDPWR.n1042 VDPWR.n1041 0.124275
R2898 VDPWR.n1060 VDPWR.n1059 0.124275
R2899 VDPWR.n1078 VDPWR.n1077 0.124275
R2900 VDPWR.n1096 VDPWR.n1095 0.124275
R2901 VDPWR.n1114 VDPWR.n1113 0.124275
R2902 VDPWR.n325 VDPWR 0.124198
R2903 VDPWR.n359 VDPWR 0.124198
R2904 VDPWR.n385 VDPWR 0.124198
R2905 VDPWR.n411 VDPWR 0.124198
R2906 VDPWR.n437 VDPWR 0.124198
R2907 VDPWR.n463 VDPWR 0.124198
R2908 VDPWR.n60 VDPWR 0.124198
R2909 VDPWR.n94 VDPWR 0.124198
R2910 VDPWR.n986 VDPWR.n973 0.121824
R2911 VDPWR.n1004 VDPWR.n969 0.121824
R2912 VDPWR.n1022 VDPWR.n965 0.121824
R2913 VDPWR.n1040 VDPWR.n961 0.121824
R2914 VDPWR.n1058 VDPWR.n957 0.121824
R2915 VDPWR.n1076 VDPWR.n953 0.121824
R2916 VDPWR.n1094 VDPWR.n949 0.121824
R2917 VDPWR.n1112 VDPWR.n945 0.121824
R2918 VDPWR.n489 VDPWR.n176 0.115083
R2919 VDPWR.n500 VDPWR.n170 0.115083
R2920 VDPWR.n128 VDPWR.n7 0.115083
R2921 VDPWR.n139 VDPWR.n1 0.115083
R2922 VDPWR VDPWR.n990 0.113245
R2923 VDPWR VDPWR.n1008 0.113245
R2924 VDPWR VDPWR.n1026 0.113245
R2925 VDPWR VDPWR.n1044 0.113245
R2926 VDPWR VDPWR.n1062 0.113245
R2927 VDPWR VDPWR.n1080 0.113245
R2928 VDPWR VDPWR.n1098 0.113245
R2929 VDPWR VDPWR.n1116 0.113245
R2930 VDPWR VDPWR.n1309 0.104667
R2931 VDPWR.n1520 VDPWR.n1519 0.10076
R2932 VDPWR.n499 VDPWR.n498 0.0899097
R2933 VDPWR.n510 VDPWR.n509 0.0899097
R2934 VDPWR.n138 VDPWR.n137 0.0899097
R2935 VDPWR.n149 VDPWR.n148 0.0899097
R2936 VDPWR.n166 VDPWR.n165 0.0826078
R2937 VDPWR.n165 VDPWR.n162 0.0777059
R2938 VDPWR.n1541 VDPWR.n1540 0.0734167
R2939 VDPWR.n1551 VDPWR.n162 0.0715784
R2940 VDPWR.n1510 VDPWR.n1509 0.0708125
R2941 VDPWR.n1504 VDPWR.n1503 0.0708125
R2942 VDPWR.n843 VDPWR 0.0708125
R2943 VDPWR VDPWR.n337 0.0695104
R2944 VDPWR.n358 VDPWR 0.0695104
R2945 VDPWR VDPWR.n371 0.0695104
R2946 VDPWR.n384 VDPWR 0.0695104
R2947 VDPWR VDPWR.n397 0.0695104
R2948 VDPWR.n410 VDPWR 0.0695104
R2949 VDPWR VDPWR.n423 0.0695104
R2950 VDPWR.n436 VDPWR 0.0695104
R2951 VDPWR VDPWR.n449 0.0695104
R2952 VDPWR.n462 VDPWR 0.0695104
R2953 VDPWR VDPWR.n475 0.0695104
R2954 VDPWR VDPWR.n72 0.0695104
R2955 VDPWR.n93 VDPWR 0.0695104
R2956 VDPWR VDPWR.n106 0.0695104
R2957 VDPWR.n1545 VDPWR.n166 0.0666765
R2958 VDPWR.n497 VDPWR.n176 0.0647361
R2959 VDPWR.n508 VDPWR.n170 0.0647361
R2960 VDPWR.n136 VDPWR.n7 0.0647361
R2961 VDPWR.n147 VDPWR.n1 0.0647361
R2962 VDPWR.n355 VDPWR 0.063
R2963 VDPWR.n124 VDPWR 0.063
R2964 VDPWR.n90 VDPWR 0.063
R2965 VDPWR.n940 VDPWR.n688 0.0577917
R2966 VDPWR.n936 VDPWR.n935 0.0577917
R2967 VDPWR.n933 VDPWR.n695 0.0577917
R2968 VDPWR.n929 VDPWR.n928 0.0577917
R2969 VDPWR.n926 VDPWR.n702 0.0577917
R2970 VDPWR.n922 VDPWR.n921 0.0577917
R2971 VDPWR.n919 VDPWR.n709 0.0577917
R2972 VDPWR.n915 VDPWR.n914 0.0577917
R2973 VDPWR.n912 VDPWR.n716 0.0577917
R2974 VDPWR.n908 VDPWR.n907 0.0577917
R2975 VDPWR.n905 VDPWR.n723 0.0577917
R2976 VDPWR.n901 VDPWR.n900 0.0577917
R2977 VDPWR.n898 VDPWR.n730 0.0577917
R2978 VDPWR.n894 VDPWR.n893 0.0577917
R2979 VDPWR.n891 VDPWR.n737 0.0577917
R2980 VDPWR.n887 VDPWR.n886 0.0577917
R2981 VDPWR.n884 VDPWR.n744 0.0577917
R2982 VDPWR.n880 VDPWR.n879 0.0577917
R2983 VDPWR.n877 VDPWR.n751 0.0577917
R2984 VDPWR.n873 VDPWR.n872 0.0577917
R2985 VDPWR.n870 VDPWR.n758 0.0577917
R2986 VDPWR.n866 VDPWR.n865 0.0577917
R2987 VDPWR.n863 VDPWR.n765 0.0577917
R2988 VDPWR.n859 VDPWR.n858 0.0577917
R2989 VDPWR.n856 VDPWR.n772 0.0577917
R2990 VDPWR.n852 VDPWR.n851 0.0577917
R2991 VDPWR.n849 VDPWR.n779 0.0577917
R2992 VDPWR.n845 VDPWR.n844 0.0577917
R2993 VDPWR.n1539 VDPWR.n1467 0.0577917
R2994 VDPWR.n1535 VDPWR.n1534 0.0577917
R2995 VDPWR.n1532 VDPWR.n1474 0.0577917
R2996 VDPWR.n1528 VDPWR.n1527 0.0577917
R2997 VDPWR.n1525 VDPWR.n1481 0.0577917
R2998 VDPWR.n1521 VDPWR.n1520 0.0577917
R2999 VDPWR.n341 VDPWR.n340 0.0577917
R3000 VDPWR.n348 VDPWR.n347 0.0577917
R3001 VDPWR.n375 VDPWR.n374 0.0577917
R3002 VDPWR.n382 VDPWR.n381 0.0577917
R3003 VDPWR.n401 VDPWR.n400 0.0577917
R3004 VDPWR.n408 VDPWR.n407 0.0577917
R3005 VDPWR.n427 VDPWR.n426 0.0577917
R3006 VDPWR.n434 VDPWR.n433 0.0577917
R3007 VDPWR.n453 VDPWR.n452 0.0577917
R3008 VDPWR.n460 VDPWR.n459 0.0577917
R3009 VDPWR.n479 VDPWR.n478 0.0577917
R3010 VDPWR.n486 VDPWR.n485 0.0577917
R3011 VDPWR.n159 VDPWR.n152 0.0577917
R3012 VDPWR.n76 VDPWR.n75 0.0577917
R3013 VDPWR.n83 VDPWR.n82 0.0577917
R3014 VDPWR.n110 VDPWR.n109 0.0577917
R3015 VDPWR.n117 VDPWR.n116 0.0577917
R3016 VDPWR.n150 VDPWR 0.0439028
R3017 VDPWR.n567 VDPWR.n550 0.0432215
R3018 VDPWR.n584 VDPWR.n545 0.0432215
R3019 VDPWR.n601 VDPWR.n540 0.0432215
R3020 VDPWR.n618 VDPWR.n535 0.0432215
R3021 VDPWR.n635 VDPWR.n530 0.0432215
R3022 VDPWR.n652 VDPWR.n525 0.0432215
R3023 VDPWR.n669 VDPWR.n520 0.0432215
R3024 VDPWR.n686 VDPWR.n515 0.0432215
R3025 VDPWR VDPWR.n488 0.0421667
R3026 VDPWR VDPWR.n127 0.0421667
R3027 VDPWR.n168 VDPWR 0.0295179
R3028 VDPWR.n1503 VDPWR.n1487 0.0278438
R3029 VDPWR.n1511 VDPWR.n1510 0.0278438
R3030 VDPWR.n1551 VDPWR 0.0201078
R3031 VDPWR.n1309 VDPWR 0.0187292
R3032 VDPWR VDPWR.n358 0.00701042
R3033 VDPWR VDPWR.n384 0.00701042
R3034 VDPWR VDPWR.n410 0.00701042
R3035 VDPWR VDPWR.n436 0.00701042
R3036 VDPWR VDPWR.n462 0.00701042
R3037 VDPWR VDPWR.n93 0.00701042
R3038 VDPWR.n160 VDPWR.n159 0.00440625
R3039 VDPWR.n987 VDPWR.n986 0.00295098
R3040 VDPWR.n1005 VDPWR.n1004 0.00295098
R3041 VDPWR.n1023 VDPWR.n1022 0.00295098
R3042 VDPWR.n1041 VDPWR.n1040 0.00295098
R3043 VDPWR.n1059 VDPWR.n1058 0.00295098
R3044 VDPWR.n1077 VDPWR.n1076 0.00295098
R3045 VDPWR.n1095 VDPWR.n1094 0.00295098
R3046 VDPWR.n1113 VDPWR.n1112 0.00295098
R3047 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 784.053
R3048 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 784.053
R3049 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 784.053
R3050 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 784.053
R3051 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 539.841
R3052 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 539.841
R3053 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 539.841
R3054 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 539.841
R3055 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 215.293
R3056 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 215.293
R3057 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 215.293
R3058 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 215.293
R3059 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 168.659
R3060 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 167.992
R3061 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 166.144
R3062 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 165.8
R3063 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 85.2499
R3064 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 85.2499
R3065 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 83.7172
R3066 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 83.7172
R3067 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 75.7282
R3068 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 66.3172
R3069 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 36.1505
R3070 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 36.1505
R3071 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 34.5438
R3072 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 34.5438
R3073 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 17.4005
R3074 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 17.4005
R3075 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 17.2391
R3076 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 9.52217
R3077 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 9.52217
R3078 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 6.39571
R3079 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 5.30824
R3080 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 4.94887
R3081 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 1.48097
R3082 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 1.06691
R3083 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.539562
R3084 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.391125
R3085 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 0.160656
R3086 tdc_0.start_buffer_0.start_buff.n11 tdc_0.start_buffer_0.start_buff.t21 543.053
R3087 tdc_0.start_buffer_0.start_buff.n12 tdc_0.start_buffer_0.start_buff.t16 543.053
R3088 tdc_0.start_buffer_0.start_buff.n10 tdc_0.start_buffer_0.start_buff.t10 543.053
R3089 tdc_0.start_buffer_0.start_buff.n1 tdc_0.start_buffer_0.start_buff.t11 539.841
R3090 tdc_0.start_buffer_0.start_buff.n0 tdc_0.start_buffer_0.start_buff.t15 539.841
R3091 tdc_0.start_buffer_0.start_buff.n4 tdc_0.start_buffer_0.start_buff.t13 539.841
R3092 tdc_0.start_buffer_0.start_buff.n3 tdc_0.start_buffer_0.start_buff.t19 539.841
R3093 tdc_0.start_buffer_0.start_buff.n11 tdc_0.start_buffer_0.start_buff.t18 221.72
R3094 tdc_0.start_buffer_0.start_buff.n12 tdc_0.start_buffer_0.start_buff.t14 221.72
R3095 tdc_0.start_buffer_0.start_buff.n10 tdc_0.start_buffer_0.start_buff.t22 221.72
R3096 tdc_0.start_buffer_0.start_buff.n13 tdc_0.start_buffer_0.start_buff.n11 218.32
R3097 tdc_0.start_buffer_0.start_buff.n13 tdc_0.start_buffer_0.start_buff.n12 217.734
R3098 tdc_0.start_buffer_0.start_buff.n1 tdc_0.start_buffer_0.start_buff.t20 215.293
R3099 tdc_0.start_buffer_0.start_buff.n0 tdc_0.start_buffer_0.start_buff.t12 215.293
R3100 tdc_0.start_buffer_0.start_buff.n4 tdc_0.start_buffer_0.start_buff.t23 215.293
R3101 tdc_0.start_buffer_0.start_buff.n3 tdc_0.start_buffer_0.start_buff.t17 215.293
R3102 tdc_0.start_buffer_0.start_buff.n14 tdc_0.start_buffer_0.start_buff.n10 213.234
R3103 tdc_0.start_buffer_0.start_buff.n6 tdc_0.start_buffer_0.start_buff.n2 166.149
R3104 tdc_0.start_buffer_0.start_buff.n6 tdc_0.start_buffer_0.start_buff.n5 165.8
R3105 tdc_0.start_buffer_0.start_buff.n18 tdc_0.start_buffer_0.start_buff.t4 85.2499
R3106 tdc_0.start_buffer_0.start_buff.n17 tdc_0.start_buffer_0.start_buff.t6 85.2499
R3107 tdc_0.start_buffer_0.start_buff.n20 tdc_0.start_buffer_0.start_buff.t7 85.2499
R3108 tdc_0.start_buffer_0.start_buff.n7 tdc_0.start_buffer_0.start_buff.t9 85.1574
R3109 tdc_0.start_buffer_0.start_buff.n9 tdc_0.start_buffer_0.start_buff.t5 83.8097
R3110 tdc_0.start_buffer_0.start_buff.n7 tdc_0.start_buffer_0.start_buff.t8 83.8097
R3111 tdc_0.start_buffer_0.start_buff.n20 tdc_0.start_buffer_0.start_buff.t3 83.7172
R3112 tdc_0.start_buffer_0.start_buff.n16 tdc_0.start_buffer_0.start_buff.t1 83.7172
R3113 tdc_0.start_buffer_0.start_buff.n18 tdc_0.start_buffer_0.start_buff.t0 83.7172
R3114 tdc_0.start_buffer_0.start_buff.n17 tdc_0.start_buffer_0.start_buff.t2 83.7172
R3115 tdc_0.start_buffer_0.start_buff.n2 tdc_0.start_buffer_0.start_buff.n1 36.1505
R3116 tdc_0.start_buffer_0.start_buff.n5 tdc_0.start_buffer_0.start_buff.n3 36.1505
R3117 tdc_0.start_buffer_0.start_buff.n2 tdc_0.start_buffer_0.start_buff.n0 34.5438
R3118 tdc_0.start_buffer_0.start_buff.n5 tdc_0.start_buffer_0.start_buff.n4 34.5438
R3119 tdc_0.start_buffer_0.start_buff.n8 tdc_0.start_buffer_0.start_buff.n6 11.8364
R3120 tdc_0.start_buffer_0.start_buff.n9 tdc_0.start_buffer_0.start_buff 8.40722
R3121 tdc_0.start_buffer_0.start_buff.n8 tdc_0.start_buffer_0.start_buff.n7 5.74235
R3122 tdc_0.start_buffer_0.start_buff.n19 tdc_0.start_buffer_0.start_buff.n17 5.16238
R3123 tdc_0.start_buffer_0.start_buff.n14 tdc_0.start_buffer_0.start_buff.n13 5.08518
R3124 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n16 4.70702
R3125 tdc_0.start_buffer_0.start_buff.n19 tdc_0.start_buffer_0.start_buff.n18 4.64452
R3126 tdc_0.start_buffer_0.start_buff.n21 tdc_0.start_buffer_0.start_buff.n20 4.64452
R3127 tdc_0.start_buffer_0.start_buff.n15 tdc_0.start_buffer_0.start_buff.n9 0.918978
R3128 tdc_0.start_buffer_0.start_buff.n21 tdc_0.start_buffer_0.start_buff.n19 0.518357
R3129 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n21 0.455857
R3130 tdc_0.start_buffer_0.start_buff.n16 tdc_0.start_buffer_0.start_buff.n15 0.3755
R3131 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n8 0.285656
R3132 tdc_0.start_buffer_0.start_buff.n15 tdc_0.start_buffer_0.start_buff.n14 0.247513
R3133 tdc_0.start_buffer_0.start_delay.n1 tdc_0.start_buffer_0.start_delay.t14 539.841
R3134 tdc_0.start_buffer_0.start_delay.n0 tdc_0.start_buffer_0.start_delay.t8 539.841
R3135 tdc_0.start_buffer_0.start_delay.n4 tdc_0.start_buffer_0.start_delay.t10 539.841
R3136 tdc_0.start_buffer_0.start_delay.n3 tdc_0.start_buffer_0.start_delay.t13 539.841
R3137 tdc_0.start_buffer_0.start_delay.n1 tdc_0.start_buffer_0.start_delay.t12 215.293
R3138 tdc_0.start_buffer_0.start_delay.n0 tdc_0.start_buffer_0.start_delay.t15 215.293
R3139 tdc_0.start_buffer_0.start_delay.n4 tdc_0.start_buffer_0.start_delay.t9 215.293
R3140 tdc_0.start_buffer_0.start_delay.n3 tdc_0.start_buffer_0.start_delay.t11 215.293
R3141 tdc_0.start_buffer_0.start_delay.n6 tdc_0.start_buffer_0.start_delay.n2 166.144
R3142 tdc_0.start_buffer_0.start_delay.n6 tdc_0.start_buffer_0.start_delay.n5 165.8
R3143 tdc_0.start_buffer_0.start_delay.n9 tdc_0.start_buffer_0.start_delay.t5 85.2499
R3144 tdc_0.start_buffer_0.start_delay.n7 tdc_0.start_buffer_0.start_delay.t6 85.2499
R3145 tdc_0.start_buffer_0.start_delay.n8 tdc_0.start_buffer_0.start_delay.t7 85.2499
R3146 tdc_0.start_buffer_0.start_delay.n11 tdc_0.start_buffer_0.start_delay.t4 84.7281
R3147 tdc_0.start_buffer_0.start_delay.n8 tdc_0.start_buffer_0.start_delay.t3 83.7172
R3148 tdc_0.start_buffer_0.start_delay.n12 tdc_0.start_buffer_0.start_delay.t0 83.7172
R3149 tdc_0.start_buffer_0.start_delay.n9 tdc_0.start_buffer_0.start_delay.t1 83.7172
R3150 tdc_0.start_buffer_0.start_delay.n7 tdc_0.start_buffer_0.start_delay.t2 83.7172
R3151 tdc_0.start_buffer_0.start_delay.n2 tdc_0.start_buffer_0.start_delay.n0 36.1505
R3152 tdc_0.start_buffer_0.start_delay.n5 tdc_0.start_buffer_0.start_delay.n3 36.1505
R3153 tdc_0.start_buffer_0.start_delay.n2 tdc_0.start_buffer_0.start_delay.n1 34.5438
R3154 tdc_0.start_buffer_0.start_delay.n5 tdc_0.start_buffer_0.start_delay.n4 34.5438
R3155 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n7 6.45821
R3156 tdc_0.start_buffer_0.start_delay.n10 tdc_0.start_buffer_0.start_delay.n8 5.16238
R3157 tdc_0.start_buffer_0.start_delay.n13 tdc_0.start_buffer_0.start_delay.n12 4.64452
R3158 tdc_0.start_buffer_0.start_delay.n10 tdc_0.start_buffer_0.start_delay.n9 4.64452
R3159 tdc_0.start_buffer_0.start_delay.n14 tdc_0.start_buffer_0.start_delay.n13 0.759429
R3160 tdc_0.start_buffer_0.start_delay.n13 tdc_0.start_buffer_0.start_delay.n10 0.518357
R3161 tdc_0.start_buffer_0.start_delay.n14 tdc_0.start_buffer_0.start_delay 0.471203
R3162 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n6 0.46925
R3163 tdc_0.start_buffer_0.start_delay.n12 tdc_0.start_buffer_0.start_delay.n11 0.3755
R3164 tdc_0.start_buffer_0.start_delay.n11 tdc_0.start_buffer_0.start_delay 0.234296
R3165 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n14 0.127453
R3166 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 628.097
R3167 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 622.766
R3168 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 523.774
R3169 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 304.647
R3170 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 304.647
R3171 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 202.44
R3172 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 169.062
R3173 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 166.237
R3174 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 84.7557
R3175 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 84.1197
R3176 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R3177 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 5.48979
R3178 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en 4.5005
R3179 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 1.09595
R3180 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 890.727
R3181 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 742.783
R3182 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 641.061
R3183 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 623.388
R3184 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 547.874
R3185 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 431.807
R3186 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 427.875
R3187 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 340.632
R3188 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 208.631
R3189 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 168.007
R3190 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R3191 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R3192 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 31.0962
R3193 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R3194 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3195 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 8.91506
R3196 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R3197 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R3198 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3199 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R3200 VGND.n1747 VGND.n166 145435
R3201 VGND.n1747 VGND.n1746 89027.6
R3202 VGND.n316 VGND.n188 35396
R3203 VGND.n1004 VGND.n166 35396
R3204 VGND.n1747 VGND.n167 31825.6
R3205 VGND.n146 VGND.n135 24188.9
R3206 VGND.n315 VGND.n137 22872.1
R3207 VGND.n1828 VGND.t30 18604.5
R3208 VGND.n168 VGND.n167 16815
R3209 VGND.n208 VGND.n188 16612
R3210 VGND.n1712 VGND.n331 14632.6
R3211 VGND.n208 VGND.t30 14477.4
R3212 VGND.n1577 VGND.t146 13628.8
R3213 VGND.n1826 VGND.t30 11061.3
R3214 VGND.n1569 VGND.n1568 9459.64
R3215 VGND.n330 VGND.n167 9082.84
R3216 VGND.n1761 VGND.t0 7799.94
R3217 VGND.n1794 VGND.n5 6289.43
R3218 VGND.n1578 VGND.n1577 6212.87
R3219 VGND.n1828 VGND.n1827 5291.8
R3220 VGND.n1577 VGND.n5 4980.04
R3221 VGND.n1709 VGND.n1578 4836.21
R3222 VGND.t155 VGND.n1828 4811.74
R3223 VGND.n314 VGND.n189 4594.02
R3224 VGND.n1569 VGND.n563 4479.04
R3225 VGND.n1570 VGND.n562 4479.04
R3226 VGND.n1571 VGND.n561 4479.04
R3227 VGND.n1572 VGND.n560 4479.04
R3228 VGND.n1573 VGND.n559 4479.04
R3229 VGND.n1574 VGND.n558 4479.04
R3230 VGND.n1575 VGND.n557 4479.04
R3231 VGND.n1576 VGND.n556 4479.04
R3232 VGND.n857 VGND.n138 4447.27
R3233 VGND.n1760 VGND.n139 4447.27
R3234 VGND.n260 VGND.n259 4447.27
R3235 VGND.n227 VGND.n226 4447.27
R3236 VGND.n1034 VGND.n520 4283.98
R3237 VGND.n1018 VGND.n520 4283.98
R3238 VGND.n696 VGND.n520 4283.98
R3239 VGND.n678 VGND.n520 4283.98
R3240 VGND.n654 VGND.n520 4283.98
R3241 VGND.n630 VGND.n520 4283.98
R3242 VGND.n606 VGND.n520 4283.98
R3243 VGND.t153 VGND.n1761 4154.59
R3244 VGND.n1548 VGND.n1163 3781.58
R3245 VGND.n1548 VGND.n1164 3781.58
R3246 VGND.n1548 VGND.n1165 3781.58
R3247 VGND.n1548 VGND.n1166 3781.58
R3248 VGND.n1548 VGND.n1167 3781.58
R3249 VGND.n1549 VGND.n1548 3781.58
R3250 VGND.n1548 VGND.n1547 3781.58
R3251 VGND.n1746 VGND.n331 3732.45
R3252 VGND.n1749 VGND.n138 3442.57
R3253 VGND.n1760 VGND.n140 3442.57
R3254 VGND.n259 VGND.n256 3442.57
R3255 VGND.n254 VGND.n227 3442.57
R3256 VGND.n1147 VGND.n563 3439.59
R3257 VGND.n331 VGND.n6 3358.06
R3258 VGND.n857 VGND.n161 3165.68
R3259 VGND.n157 VGND.n139 3165.68
R3260 VGND.n260 VGND.n220 3165.68
R3261 VGND.n230 VGND.n226 3165.68
R3262 VGND.n1161 VGND.n563 3093.4
R3263 VGND.n1470 VGND.n562 3093.4
R3264 VGND.n1458 VGND.n561 3093.4
R3265 VGND.n1446 VGND.n560 3093.4
R3266 VGND.n1434 VGND.n559 3093.4
R3267 VGND.n1422 VGND.n558 3093.4
R3268 VGND.n1409 VGND.n557 3093.4
R3269 VGND.n1535 VGND.n556 3093.4
R3270 VGND.n1236 VGND.n521 3089.56
R3271 VGND.n1386 VGND.n527 3089.56
R3272 VGND.n1376 VGND.n522 3089.56
R3273 VGND.n1351 VGND.n526 3089.56
R3274 VGND.n1326 VGND.n523 3089.56
R3275 VGND.n1301 VGND.n525 3089.56
R3276 VGND.n1727 VGND.n519 3089.56
R3277 VGND.n1725 VGND.n529 3089.56
R3278 VGND.n1235 VGND.n1170 2843.1
R3279 VGND.n1385 VGND.n1171 2843.1
R3280 VGND.n1375 VGND.n1172 2843.1
R3281 VGND.n1350 VGND.n1173 2843.1
R3282 VGND.n1325 VGND.n1174 2843.1
R3283 VGND.n1300 VGND.n1175 2843.1
R3284 VGND.n1177 VGND.n1176 2843.1
R3285 VGND.n1169 VGND.n536 2843.1
R3286 VGND.n1827 VGND.n1826 2773.54
R3287 VGND.n1711 VGND.n1710 2755.48
R3288 VGND.n1568 VGND.n565 2713.47
R3289 VGND.n314 VGND.n313 2502.61
R3290 VGND.n331 VGND.n330 2480.88
R3291 VGND.n1568 VGND.n1567 2378.68
R3292 VGND.n1240 VGND.n521 2350.81
R3293 VGND.n1226 VGND.n527 2350.81
R3294 VGND.n1365 VGND.n522 2350.81
R3295 VGND.n1340 VGND.n526 2350.81
R3296 VGND.n1315 VGND.n523 2350.81
R3297 VGND.n1290 VGND.n525 2350.81
R3298 VGND.n1727 VGND.n518 2350.81
R3299 VGND.n1725 VGND.n528 2350.81
R3300 VGND.n1749 VGND.n162 2206.4
R3301 VGND.n158 VGND.n140 2206.4
R3302 VGND.n256 VGND.n223 2206.4
R3303 VGND.n254 VGND.n225 2206.4
R3304 VGND.n238 VGND.n136 2152.16
R3305 VGND.n151 VGND.n146 2067.34
R3306 VGND.n1600 VGND.n1595 2058.56
R3307 VGND.n1693 VGND.n1595 2058.56
R3308 VGND.n1690 VGND.n1603 2058.56
R3309 VGND.n1622 VGND.n1603 2058.56
R3310 VGND.n1624 VGND.n1619 2058.56
R3311 VGND.n1675 VGND.n1619 2058.56
R3312 VGND.n1672 VGND.n1627 2058.56
R3313 VGND.n1649 VGND.n1627 2058.56
R3314 VGND.n1651 VGND.n1646 2058.56
R3315 VGND.n1657 VGND.n1646 2058.56
R3316 VGND.n1792 VGND.n75 2058.56
R3317 VGND.n1654 VGND.n75 2058.56
R3318 VGND.n1598 VGND.n1579 2058.56
R3319 VGND.n1707 VGND.n1579 2058.56
R3320 VGND.n1566 VGND.n566 2058.56
R3321 VGND.n1148 VGND.n566 2058.56
R3322 VGND.n1160 VGND.n1159 2058.56
R3323 VGND.n1551 VGND.n1159 2058.56
R3324 VGND.n1471 VGND.n1466 2058.56
R3325 VGND.n1467 VGND.n1466 2058.56
R3326 VGND.n1459 VGND.n1454 2058.56
R3327 VGND.n1455 VGND.n1454 2058.56
R3328 VGND.n1447 VGND.n1442 2058.56
R3329 VGND.n1443 VGND.n1442 2058.56
R3330 VGND.n1435 VGND.n1430 2058.56
R3331 VGND.n1431 VGND.n1430 2058.56
R3332 VGND.n1423 VGND.n1418 2058.56
R3333 VGND.n1419 VGND.n1418 2058.56
R3334 VGND.n1410 VGND.n1401 2058.56
R3335 VGND.n1545 VGND.n1401 2058.56
R3336 VGND.n1533 VGND.n1532 2058.56
R3337 VGND.n1534 VGND.n1533 2058.56
R3338 VGND.n1189 VGND.n1188 2029.1
R3339 VGND.n1393 VGND.n1220 2029.1
R3340 VGND.n1192 VGND.n1191 2029.1
R3341 VGND.n1218 VGND.n1217 2029.1
R3342 VGND.n1195 VGND.n1194 2029.1
R3343 VGND.n1215 VGND.n1214 2029.1
R3344 VGND.n1212 VGND.n1197 2029.1
R3345 VGND.n1395 VGND.n1186 2029.1
R3346 VGND.n1251 VGND.n1184 1929.2
R3347 VGND.n1230 VGND.n1183 1929.2
R3348 VGND.n1366 VGND.n1182 1929.2
R3349 VGND.n1341 VGND.n1181 1929.2
R3350 VGND.n1316 VGND.n1180 1929.2
R3351 VGND.n1291 VGND.n1179 1929.2
R3352 VGND.n1204 VGND.n1178 1929.2
R3353 VGND.n1399 VGND.n1185 1929.2
R3354 VGND.n509 VGND.n6 1814.76
R3355 VGND.n1549 VGND.n562 1809.14
R3356 VGND.n1167 VGND.n561 1809.14
R3357 VGND.n1166 VGND.n560 1809.14
R3358 VGND.n1165 VGND.n559 1809.14
R3359 VGND.n1164 VGND.n558 1809.14
R3360 VGND.n1163 VGND.n557 1809.14
R3361 VGND.n1547 VGND.n556 1809.14
R3362 VGND.n1568 VGND.n564 1741.86
R3363 VGND.n1189 VGND.n1187 1718.82
R3364 VGND.n1393 VGND.n1219 1718.82
R3365 VGND.n1192 VGND.n1190 1718.82
R3366 VGND.n1218 VGND.n1216 1718.82
R3367 VGND.n1195 VGND.n1193 1718.82
R3368 VGND.n1215 VGND.n1213 1718.82
R3369 VGND.n1212 VGND.n1196 1718.82
R3370 VGND.n1395 VGND.n535 1718.82
R3371 VGND.n1763 VGND.n135 1708.68
R3372 VGND.n1829 VGND.n3 1707.33
R3373 VGND.n1831 VGND.n3 1707.33
R3374 VGND.n1764 VGND.n133 1707.33
R3375 VGND.n1764 VGND.n134 1707.33
R3376 VGND.n188 VGND.n6 1644.04
R3377 VGND.n1550 VGND.n1549 1630.46
R3378 VGND.n1468 VGND.n1167 1630.46
R3379 VGND.n1456 VGND.n1166 1630.46
R3380 VGND.n1444 VGND.n1165 1630.46
R3381 VGND.n1432 VGND.n1164 1630.46
R3382 VGND.n1420 VGND.n1163 1630.46
R3383 VGND.n1547 VGND.n1546 1630.46
R3384 VGND.n185 VGND.n180 1626.7
R3385 VGND.n318 VGND.n180 1626.7
R3386 VGND.n312 VGND.n192 1626.7
R3387 VGND.n312 VGND.n193 1626.7
R3388 VGND.n302 VGND.n190 1626.7
R3389 VGND.n304 VGND.n190 1626.7
R3390 VGND.n1000 VGND.n737 1626.7
R3391 VGND.n1006 VGND.n737 1626.7
R3392 VGND.n975 VGND.n770 1626.7
R3393 VGND.n977 VGND.n770 1626.7
R3394 VGND.n974 VGND.n790 1626.7
R3395 VGND.n790 VGND.n772 1626.7
R3396 VGND.n953 VGND.n789 1626.7
R3397 VGND.n953 VGND.n773 1626.7
R3398 VGND.n808 VGND.n788 1626.7
R3399 VGND.n808 VGND.n774 1626.7
R3400 VGND.n931 VGND.n787 1626.7
R3401 VGND.n931 VGND.n775 1626.7
R3402 VGND.n822 VGND.n786 1626.7
R3403 VGND.n822 VGND.n776 1626.7
R3404 VGND.n909 VGND.n785 1626.7
R3405 VGND.n909 VGND.n777 1626.7
R3406 VGND.n836 VGND.n784 1626.7
R3407 VGND.n836 VGND.n778 1626.7
R3408 VGND.n887 VGND.n783 1626.7
R3409 VGND.n887 VGND.n779 1626.7
R3410 VGND.n850 VGND.n782 1626.7
R3411 VGND.n850 VGND.n780 1626.7
R3412 VGND.n1016 VGND.n726 1626.7
R3413 VGND.n998 VGND.n726 1626.7
R3414 VGND.n328 VGND.n169 1626.7
R3415 VGND.n183 VGND.n169 1626.7
R3416 VGND.n1761 VGND.n136 1617.44
R3417 VGND.n1253 VGND.n1240 1562.99
R3418 VGND.n1232 VGND.n1226 1562.99
R3419 VGND.n1368 VGND.n1365 1562.99
R3420 VGND.n1343 VGND.n1340 1562.99
R3421 VGND.n1318 VGND.n1315 1562.99
R3422 VGND.n1293 VGND.n1290 1562.99
R3423 VGND.n1202 VGND.n518 1562.99
R3424 VGND.n1714 VGND.n528 1562.99
R3425 VGND.n1570 VGND.n1569 1482.26
R3426 VGND.n1571 VGND.n1570 1482.26
R3427 VGND.n1572 VGND.n1571 1482.26
R3428 VGND.n1573 VGND.n1572 1482.26
R3429 VGND.n1574 VGND.n1573 1482.26
R3430 VGND.n1575 VGND.n1574 1482.26
R3431 VGND.n1576 VGND.n1575 1482.26
R3432 VGND.n1578 VGND.n1576 1458.22
R3433 VGND.n1753 VGND.n162 1438.1
R3434 VGND.n1755 VGND.n158 1438.1
R3435 VGND.n264 VGND.n223 1438.1
R3436 VGND.n225 VGND.n224 1438.1
R3437 VGND.n1793 VGND.n1791 1396.01
R3438 VGND.n1825 VGND.n1824 1325.13
R3439 VGND.n1710 VGND.n555 1263.93
R3440 VGND.n1709 VGND.n1708 1228.29
R3441 VGND.n1188 VGND.n1184 1210.97
R3442 VGND.n1220 VGND.n1183 1210.97
R3443 VGND.n1191 VGND.n1182 1210.97
R3444 VGND.n1217 VGND.n1181 1210.97
R3445 VGND.n1194 VGND.n1180 1210.97
R3446 VGND.n1214 VGND.n1179 1210.97
R3447 VGND.n1197 VGND.n1178 1210.97
R3448 VGND.n1399 VGND.n1186 1210.97
R3449 VGND.n1188 VGND.n1170 1199.38
R3450 VGND.n1220 VGND.n1171 1199.38
R3451 VGND.n1191 VGND.n1172 1199.38
R3452 VGND.n1217 VGND.n1173 1199.38
R3453 VGND.n1194 VGND.n1174 1199.38
R3454 VGND.n1214 VGND.n1175 1199.38
R3455 VGND.n1197 VGND.n1177 1199.38
R3456 VGND.n1186 VGND.n1169 1199.38
R3457 VGND.n1827 VGND.n5 1074.72
R3458 VGND.n1753 VGND.n161 1065.44
R3459 VGND.n1755 VGND.n157 1065.44
R3460 VGND.n264 VGND.n220 1065.44
R3461 VGND.n230 VGND.n224 1065.44
R3462 VGND.n300 VGND.n283 1058.19
R3463 VGND.n283 VGND.n204 1058.19
R3464 VGND.n288 VGND.n282 1058.19
R3465 VGND.n288 VGND.n205 1058.19
R3466 VGND.n281 VGND.n210 1058.19
R3467 VGND.n210 VGND.n206 1058.19
R3468 VGND.n215 VGND.n209 1058.19
R3469 VGND.n215 VGND.n207 1058.19
R3470 VGND.n240 VGND.n237 1058.19
R3471 VGND.n242 VGND.n237 1058.19
R3472 VGND.n152 VGND.n145 1058.19
R3473 VGND.n150 VGND.n145 1058.19
R3474 VGND.n989 VGND.n740 1058.19
R3475 VGND.n991 VGND.n740 1058.19
R3476 VGND.n988 VGND.n763 1058.19
R3477 VGND.n763 VGND.n742 1058.19
R3478 VGND.n797 VGND.n762 1058.19
R3479 VGND.n797 VGND.n743 1058.19
R3480 VGND.n800 VGND.n761 1058.19
R3481 VGND.n800 VGND.n744 1058.19
R3482 VGND.n811 VGND.n760 1058.19
R3483 VGND.n811 VGND.n745 1058.19
R3484 VGND.n814 VGND.n759 1058.19
R3485 VGND.n814 VGND.n746 1058.19
R3486 VGND.n825 VGND.n758 1058.19
R3487 VGND.n825 VGND.n747 1058.19
R3488 VGND.n828 VGND.n757 1058.19
R3489 VGND.n828 VGND.n748 1058.19
R3490 VGND.n839 VGND.n756 1058.19
R3491 VGND.n839 VGND.n749 1058.19
R3492 VGND.n842 VGND.n755 1058.19
R3493 VGND.n842 VGND.n750 1058.19
R3494 VGND.n853 VGND.n754 1058.19
R3495 VGND.n853 VGND.n751 1058.19
R3496 VGND.n856 VGND.n753 1058.19
R3497 VGND.n856 VGND.n752 1058.19
R3498 VGND.n1804 VGND.n12 1058.19
R3499 VGND.n510 VGND.n343 1058.19
R3500 VGND.n1773 VGND.n79 1058.19
R3501 VGND.n1790 VGND.n84 1058.19
R3502 VGND.n1826 VGND.n1825 987.279
R3503 VGND.n1567 VGND.t343 815.229
R3504 VGND.n1146 VGND.t414 815.229
R3505 VGND.t530 VGND.n1146 815.229
R3506 VGND.n1147 VGND.t281 815.229
R3507 VGND.t520 VGND.n1161 815.229
R3508 VGND.n1162 VGND.t518 815.229
R3509 VGND.t540 VGND.n1162 815.229
R3510 VGND.n1550 VGND.t309 815.229
R3511 VGND.n1470 VGND.t181 815.229
R3512 VGND.t183 VGND.n1469 815.229
R3513 VGND.n1469 VGND.t433 815.229
R3514 VGND.t233 VGND.n1468 815.229
R3515 VGND.n1458 VGND.t89 815.229
R3516 VGND.t316 VGND.n1457 815.229
R3517 VGND.n1457 VGND.t461 815.229
R3518 VGND.t421 VGND.n1456 815.229
R3519 VGND.n1446 VGND.t50 815.229
R3520 VGND.t258 VGND.n1445 815.229
R3521 VGND.n1445 VGND.t391 815.229
R3522 VGND.t389 VGND.n1444 815.229
R3523 VGND.n1434 VGND.t262 815.229
R3524 VGND.t268 VGND.n1433 815.229
R3525 VGND.n1433 VGND.t219 815.229
R3526 VGND.t508 VGND.n1432 815.229
R3527 VGND.n1422 VGND.t64 815.229
R3528 VGND.t77 VGND.n1421 815.229
R3529 VGND.n1421 VGND.t514 815.229
R3530 VGND.t516 VGND.n1420 815.229
R3531 VGND.n1409 VGND.t213 815.229
R3532 VGND.t217 VGND.n1408 815.229
R3533 VGND.n1408 VGND.t488 815.229
R3534 VGND.n1546 VGND.t58 815.229
R3535 VGND.t9 VGND.n1535 815.229
R3536 VGND.n1536 VGND.t11 815.229
R3537 VGND.n1536 VGND.t62 815.229
R3538 VGND.n62 VGND.n61 760.639
R3539 VGND.n56 VGND.n55 760.639
R3540 VGND.n50 VGND.n49 760.639
R3541 VGND.n44 VGND.n43 760.639
R3542 VGND.n38 VGND.n37 760.639
R3543 VGND.n32 VGND.n31 760.639
R3544 VGND.n26 VGND.n25 760.639
R3545 VGND.n470 VGND.n16 760.639
R3546 VGND.n466 VGND.n465 760.639
R3547 VGND.n460 VGND.n459 760.639
R3548 VGND.n454 VGND.n453 760.639
R3549 VGND.n448 VGND.n447 760.639
R3550 VGND.n442 VGND.n441 760.639
R3551 VGND.n436 VGND.n435 760.639
R3552 VGND.n430 VGND.n429 760.639
R3553 VGND.n424 VGND.n423 760.639
R3554 VGND.n418 VGND.n417 760.639
R3555 VGND.n412 VGND.n411 760.639
R3556 VGND.n406 VGND.n405 760.639
R3557 VGND.n400 VGND.n399 760.639
R3558 VGND.n394 VGND.n393 760.639
R3559 VGND.n388 VGND.n387 760.639
R3560 VGND.n382 VGND.n381 760.639
R3561 VGND.n376 VGND.n364 760.639
R3562 VGND.n366 VGND.n363 760.639
R3563 VGND.n368 VGND.n344 760.639
R3564 VGND.n20 VGND.n17 760.639
R3565 VGND.n124 VGND.n123 760.639
R3566 VGND.n118 VGND.n117 760.639
R3567 VGND.n112 VGND.n111 760.639
R3568 VGND.n106 VGND.n105 760.639
R3569 VGND.n100 VGND.n99 760.639
R3570 VGND.n94 VGND.n93 760.639
R3571 VGND.n88 VGND.n85 760.639
R3572 VGND.n1050 VGND.n712 744.222
R3573 VGND.n1025 VGND.n711 744.222
R3574 VGND.n1022 VGND.n713 744.222
R3575 VGND.n334 VGND.n333 744.222
R3576 VGND.n1738 VGND.n337 744.222
R3577 VGND.n1042 VGND.n1033 744.222
R3578 VGND.n1128 VGND.n581 744.222
R3579 VGND.n589 VGND.n580 744.222
R3580 VGND.n586 VGND.n583 744.222
R3581 VGND.n1115 VGND.n603 744.222
R3582 VGND.n613 VGND.n602 744.222
R3583 VGND.n610 VGND.n604 744.222
R3584 VGND.n1102 VGND.n627 744.222
R3585 VGND.n637 VGND.n626 744.222
R3586 VGND.n634 VGND.n628 744.222
R3587 VGND.n1089 VGND.n651 744.222
R3588 VGND.n661 VGND.n650 744.222
R3589 VGND.n658 VGND.n652 744.222
R3590 VGND.n1076 VGND.n675 744.222
R3591 VGND.n685 VGND.n674 744.222
R3592 VGND.n682 VGND.n676 744.222
R3593 VGND.n717 VGND.n716 744.222
R3594 VGND.n718 VGND.n699 744.222
R3595 VGND.n1071 VGND.n695 744.222
R3596 VGND.n1252 VGND.n1251 742.855
R3597 VGND.n1231 VGND.n1230 742.855
R3598 VGND.n1367 VGND.n1366 742.855
R3599 VGND.n1342 VGND.n1341 742.855
R3600 VGND.n1317 VGND.n1316 742.855
R3601 VGND.n1292 VGND.n1291 742.855
R3602 VGND.n1204 VGND.n1203 742.855
R3603 VGND.n1185 VGND.n553 742.855
R3604 VGND.n1252 VGND.n552 719.461
R3605 VGND.n1231 VGND.n551 719.461
R3606 VGND.n1367 VGND.n550 719.461
R3607 VGND.n1342 VGND.n549 719.461
R3608 VGND.n1317 VGND.n548 719.461
R3609 VGND.n1292 VGND.n547 719.461
R3610 VGND.n1203 VGND.n546 719.461
R3611 VGND.n1718 VGND.n553 719.461
R3612 VGND.n1601 VGND.n1599 631.795
R3613 VGND.n1692 VGND.n1691 631.795
R3614 VGND.n1625 VGND.n1623 631.795
R3615 VGND.n1674 VGND.n1673 631.795
R3616 VGND.n1652 VGND.n1650 631.795
R3617 VGND.n1656 VGND.n1655 631.795
R3618 VGND.n728 VGND.t562 607.409
R3619 VGND.n171 VGND.t563 607.409
R3620 VGND.n1035 VGND.n1032 587.761
R3621 VGND.n1744 VGND.n1743 587.761
R3622 VGND.n1021 VGND.n714 587.761
R3623 VGND.n1027 VGND.n710 587.761
R3624 VGND.n681 VGND.n677 587.761
R3625 VGND.n687 VGND.n673 587.761
R3626 VGND.n657 VGND.n653 587.761
R3627 VGND.n663 VGND.n649 587.761
R3628 VGND.n633 VGND.n629 587.761
R3629 VGND.n639 VGND.n625 587.761
R3630 VGND.n609 VGND.n605 587.761
R3631 VGND.n615 VGND.n601 587.761
R3632 VGND.n585 VGND.n584 587.761
R3633 VGND.n591 VGND.n579 587.761
R3634 VGND.n697 VGND.n694 587.761
R3635 VGND.n724 VGND.n723 587.761
R3636 VGND.n725 VGND.n724 585
R3637 VGND.n698 VGND.n697 585
R3638 VGND.n688 VGND.n687 585
R3639 VGND.n681 VGND.n680 585
R3640 VGND.n664 VGND.n663 585
R3641 VGND.n657 VGND.n656 585
R3642 VGND.n640 VGND.n639 585
R3643 VGND.n633 VGND.n632 585
R3644 VGND.n616 VGND.n615 585
R3645 VGND.n609 VGND.n608 585
R3646 VGND.n592 VGND.n591 585
R3647 VGND.n585 VGND.n564 585
R3648 VGND.n1745 VGND.n1744 585
R3649 VGND.n1036 VGND.n1035 585
R3650 VGND.n1028 VGND.n1027 585
R3651 VGND.n1021 VGND.n1020 585
R3652 VGND.n1235 VGND.n538 561.451
R3653 VGND.n1385 VGND.n539 561.451
R3654 VGND.n1375 VGND.n540 561.451
R3655 VGND.n1350 VGND.n541 561.451
R3656 VGND.n1325 VGND.n542 561.451
R3657 VGND.n1300 VGND.n543 561.451
R3658 VGND.n1176 VGND.n544 561.451
R3659 VGND.n1720 VGND.n536 561.451
R3660 VGND.n1597 VGND.t272 549.061
R3661 VGND.t172 VGND.n1597 549.061
R3662 VGND.n1599 VGND.t535 549.061
R3663 VGND.t247 VGND.n1601 549.061
R3664 VGND.n1602 VGND.t249 549.061
R3665 VGND.t70 VGND.n1602 549.061
R3666 VGND.n1692 VGND.t215 549.061
R3667 VGND.n1691 VGND.t306 549.061
R3668 VGND.n1621 VGND.t427 549.061
R3669 VGND.t141 VGND.n1621 549.061
R3670 VGND.n1623 VGND.t506 549.061
R3671 VGND.t178 VGND.n1625 549.061
R3672 VGND.n1626 VGND.t101 549.061
R3673 VGND.t278 VGND.n1626 549.061
R3674 VGND.n1674 VGND.t332 549.061
R3675 VGND.n1673 VGND.t251 549.061
R3676 VGND.n1648 VGND.t544 549.061
R3677 VGND.t56 VGND.n1648 549.061
R3678 VGND.n1650 VGND.t454 549.061
R3679 VGND.t121 VGND.n1652 549.061
R3680 VGND.n1653 VGND.t68 549.061
R3681 VGND.t328 VGND.n1653 549.061
R3682 VGND.n1656 VGND.t330 549.061
R3683 VGND.n1655 VGND.t383 549.061
R3684 VGND.n1795 VGND.t374 549.061
R3685 VGND.n1795 VGND.t366 549.061
R3686 VGND.n1187 VGND.n552 541.75
R3687 VGND.n1219 VGND.n551 541.75
R3688 VGND.n1190 VGND.n550 541.75
R3689 VGND.n1216 VGND.n549 541.75
R3690 VGND.n1193 VGND.n548 541.75
R3691 VGND.n1213 VGND.n547 541.75
R3692 VGND.n1196 VGND.n546 541.75
R3693 VGND.n1718 VGND.n535 541.75
R3694 VGND.n1023 VGND.n1022 540.784
R3695 VGND.n1023 VGND.n711 540.784
R3696 VGND.n1039 VGND.n1033 540.784
R3697 VGND.n1039 VGND.n337 540.784
R3698 VGND.n587 VGND.n586 540.784
R3699 VGND.n587 VGND.n580 540.784
R3700 VGND.n611 VGND.n610 540.784
R3701 VGND.n611 VGND.n602 540.784
R3702 VGND.n635 VGND.n634 540.784
R3703 VGND.n635 VGND.n626 540.784
R3704 VGND.n659 VGND.n658 540.784
R3705 VGND.n659 VGND.n650 540.784
R3706 VGND.n683 VGND.n682 540.784
R3707 VGND.n683 VGND.n674 540.784
R3708 VGND.n1068 VGND.n695 540.784
R3709 VGND.n1068 VGND.n699 540.784
R3710 VGND.n1053 VGND.n711 534.99
R3711 VGND.n1053 VGND.n712 534.99
R3712 VGND.n1741 VGND.n337 534.99
R3713 VGND.n1741 VGND.n333 534.99
R3714 VGND.n1131 VGND.n580 534.99
R3715 VGND.n1131 VGND.n581 534.99
R3716 VGND.n1118 VGND.n602 534.99
R3717 VGND.n1118 VGND.n603 534.99
R3718 VGND.n1105 VGND.n626 534.99
R3719 VGND.n1105 VGND.n627 534.99
R3720 VGND.n1092 VGND.n650 534.99
R3721 VGND.n1092 VGND.n651 534.99
R3722 VGND.n1079 VGND.n674 534.99
R3723 VGND.n1079 VGND.n675 534.99
R3724 VGND.n721 VGND.n699 534.99
R3725 VGND.n721 VGND.n717 534.99
R3726 VGND.n1187 VGND.n538 507.276
R3727 VGND.n1219 VGND.n539 507.276
R3728 VGND.n1190 VGND.n540 507.276
R3729 VGND.n1216 VGND.n541 507.276
R3730 VGND.n1193 VGND.n542 507.276
R3731 VGND.n1213 VGND.n543 507.276
R3732 VGND.n1196 VGND.n544 507.276
R3733 VGND.n1720 VGND.n535 507.276
R3734 VGND.t288 VGND.t343 491.372
R3735 VGND.t211 VGND.t288 491.372
R3736 VGND.t414 VGND.t211 491.372
R3737 VGND.t44 VGND.t530 491.372
R3738 VGND.t164 VGND.t44 491.372
R3739 VGND.t281 VGND.t164 491.372
R3740 VGND.t522 VGND.t520 491.372
R3741 VGND.t60 VGND.t522 491.372
R3742 VGND.t518 VGND.t60 491.372
R3743 VGND.t538 VGND.t540 491.372
R3744 VGND.t312 VGND.t538 491.372
R3745 VGND.t309 VGND.t312 491.372
R3746 VGND.t181 VGND.t323 491.372
R3747 VGND.t323 VGND.t52 491.372
R3748 VGND.t52 VGND.t183 491.372
R3749 VGND.t433 VGND.t449 491.372
R3750 VGND.t449 VGND.t447 491.372
R3751 VGND.t447 VGND.t233 491.372
R3752 VGND.t89 VGND.t314 491.372
R3753 VGND.t314 VGND.t72 491.372
R3754 VGND.t72 VGND.t316 491.372
R3755 VGND.t461 VGND.t84 491.372
R3756 VGND.t84 VGND.t423 491.372
R3757 VGND.t423 VGND.t421 491.372
R3758 VGND.t50 VGND.t352 491.372
R3759 VGND.t352 VGND.t176 491.372
R3760 VGND.t176 VGND.t258 491.372
R3761 VGND.t391 VGND.t385 491.372
R3762 VGND.t385 VGND.t387 491.372
R3763 VGND.t387 VGND.t389 491.372
R3764 VGND.t262 VGND.t264 491.372
R3765 VGND.t264 VGND.t266 491.372
R3766 VGND.t266 VGND.t268 491.372
R3767 VGND.t219 VGND.t510 491.372
R3768 VGND.t510 VGND.t350 491.372
R3769 VGND.t350 VGND.t508 491.372
R3770 VGND.t64 VGND.t110 491.372
R3771 VGND.t110 VGND.t79 491.372
R3772 VGND.t79 VGND.t77 491.372
R3773 VGND.t514 VGND.t486 491.372
R3774 VGND.t486 VGND.t39 491.372
R3775 VGND.t39 VGND.t516 491.372
R3776 VGND.t213 VGND.t48 491.372
R3777 VGND.t48 VGND.t239 491.372
R3778 VGND.t239 VGND.t217 491.372
R3779 VGND.t488 VGND.t468 491.372
R3780 VGND.t468 VGND.t54 491.372
R3781 VGND.t54 VGND.t58 491.372
R3782 VGND.t19 VGND.t9 491.372
R3783 VGND.t5 VGND.t19 491.372
R3784 VGND.t11 VGND.t5 491.372
R3785 VGND.t62 VGND.t81 471.786
R3786 VGND.n314 VGND.n136 455.522
R3787 VGND.n1003 VGND.n159 442.918
R3788 VGND.n263 VGND.n189 430.216
R3789 VGND.n259 VGND.t30 377.098
R3790 VGND.n227 VGND.t30 377.098
R3791 VGND.n1253 VGND.n1252 356.277
R3792 VGND.n1232 VGND.n1231 356.277
R3793 VGND.n1368 VGND.n1367 356.277
R3794 VGND.n1343 VGND.n1342 356.277
R3795 VGND.n1318 VGND.n1317 356.277
R3796 VGND.n1293 VGND.n1292 356.277
R3797 VGND.n1203 VGND.n1202 356.277
R3798 VGND.n1714 VGND.n553 356.277
R3799 VGND.t188 VGND.n555 346.868
R3800 VGND.n1708 VGND.t270 346.868
R3801 VGND.n261 VGND.n255 334.05
R3802 VGND.t272 VGND.t21 330.94
R3803 VGND.t463 VGND.t172 330.94
R3804 VGND.t205 VGND.t463 330.94
R3805 VGND.t535 VGND.t205 330.94
R3806 VGND.t66 VGND.t247 330.94
R3807 VGND.t231 VGND.t66 330.94
R3808 VGND.t249 VGND.t231 330.94
R3809 VGND.t108 VGND.t70 330.94
R3810 VGND.t500 VGND.t108 330.94
R3811 VGND.t215 VGND.t500 330.94
R3812 VGND.t419 VGND.t306 330.94
R3813 VGND.t304 VGND.t419 330.94
R3814 VGND.t427 VGND.t304 330.94
R3815 VGND.t138 VGND.t141 330.94
R3816 VGND.t112 VGND.t138 330.94
R3817 VGND.t506 VGND.t112 330.94
R3818 VGND.t103 VGND.t178 330.94
R3819 VGND.t196 VGND.t103 330.94
R3820 VGND.t101 VGND.t196 330.94
R3821 VGND.t431 VGND.t278 330.94
R3822 VGND.t429 VGND.t431 330.94
R3823 VGND.t332 VGND.t429 330.94
R3824 VGND.t300 VGND.t251 330.94
R3825 VGND.t254 VGND.t300 330.94
R3826 VGND.t544 VGND.t254 330.94
R3827 VGND.t479 VGND.t56 330.94
R3828 VGND.t321 VGND.t479 330.94
R3829 VGND.t454 VGND.t321 330.94
R3830 VGND.t318 VGND.t121 330.94
R3831 VGND.t46 VGND.t318 330.94
R3832 VGND.t68 VGND.t46 330.94
R3833 VGND.t276 VGND.t328 330.94
R3834 VGND.t274 VGND.t276 330.94
R3835 VGND.t330 VGND.t274 330.94
R3836 VGND.t383 VGND.t377 330.94
R3837 VGND.t377 VGND.t380 330.94
R3838 VGND.t380 VGND.t374 330.94
R3839 VGND.t366 VGND.t368 330.94
R3840 VGND.t0 VGND.n138 325.082
R3841 VGND.t0 VGND.n1760 325.082
R3842 VGND.n728 VGND.t17 321.423
R3843 VGND.n171 VGND.t15 321.423
R3844 VGND.n1791 VGND.n80 303.616
R3845 VGND.n510 VGND.n344 297.553
R3846 VGND.n345 VGND.n344 297.553
R3847 VGND.n363 VGND.n345 297.553
R3848 VGND.n508 VGND.n363 297.553
R3849 VGND.n508 VGND.n364 297.553
R3850 VGND.n364 VGND.n346 297.553
R3851 VGND.n381 VGND.n346 297.553
R3852 VGND.n381 VGND.n362 297.553
R3853 VGND.n387 VGND.n362 297.553
R3854 VGND.n387 VGND.n347 297.553
R3855 VGND.n393 VGND.n347 297.553
R3856 VGND.n393 VGND.n361 297.553
R3857 VGND.n399 VGND.n361 297.553
R3858 VGND.n399 VGND.n348 297.553
R3859 VGND.n405 VGND.n348 297.553
R3860 VGND.n405 VGND.n360 297.553
R3861 VGND.n411 VGND.n360 297.553
R3862 VGND.n411 VGND.n349 297.553
R3863 VGND.n417 VGND.n349 297.553
R3864 VGND.n417 VGND.n359 297.553
R3865 VGND.n423 VGND.n359 297.553
R3866 VGND.n423 VGND.n350 297.553
R3867 VGND.n429 VGND.n350 297.553
R3868 VGND.n429 VGND.n358 297.553
R3869 VGND.n435 VGND.n358 297.553
R3870 VGND.n435 VGND.n351 297.553
R3871 VGND.n441 VGND.n351 297.553
R3872 VGND.n441 VGND.n357 297.553
R3873 VGND.n447 VGND.n357 297.553
R3874 VGND.n447 VGND.n352 297.553
R3875 VGND.n453 VGND.n352 297.553
R3876 VGND.n453 VGND.n356 297.553
R3877 VGND.n459 VGND.n356 297.553
R3878 VGND.n459 VGND.n353 297.553
R3879 VGND.n465 VGND.n353 297.553
R3880 VGND.n465 VGND.n355 297.553
R3881 VGND.n355 VGND.n16 297.553
R3882 VGND.n1823 VGND.n16 297.553
R3883 VGND.n1823 VGND.n17 297.553
R3884 VGND.n17 VGND.n7 297.553
R3885 VGND.n25 VGND.n7 297.553
R3886 VGND.n25 VGND.n15 297.553
R3887 VGND.n31 VGND.n15 297.553
R3888 VGND.n31 VGND.n8 297.553
R3889 VGND.n37 VGND.n8 297.553
R3890 VGND.n37 VGND.n14 297.553
R3891 VGND.n43 VGND.n14 297.553
R3892 VGND.n43 VGND.n9 297.553
R3893 VGND.n49 VGND.n9 297.553
R3894 VGND.n49 VGND.n13 297.553
R3895 VGND.n55 VGND.n13 297.553
R3896 VGND.n55 VGND.n10 297.553
R3897 VGND.n61 VGND.n10 297.553
R3898 VGND.n61 VGND.n12 297.553
R3899 VGND.n1790 VGND.n85 297.553
R3900 VGND.n85 VGND.n76 297.553
R3901 VGND.n93 VGND.n76 297.553
R3902 VGND.n93 VGND.n83 297.553
R3903 VGND.n99 VGND.n83 297.553
R3904 VGND.n99 VGND.n77 297.553
R3905 VGND.n105 VGND.n77 297.553
R3906 VGND.n105 VGND.n82 297.553
R3907 VGND.n111 VGND.n82 297.553
R3908 VGND.n111 VGND.n78 297.553
R3909 VGND.n117 VGND.n78 297.553
R3910 VGND.n117 VGND.n81 297.553
R3911 VGND.n123 VGND.n81 297.553
R3912 VGND.n123 VGND.n79 297.553
R3913 VGND.n158 VGND.n142 292.5
R3914 VGND.n771 VGND.n158 292.5
R3915 VGND.n1751 VGND.n162 292.5
R3916 VGND.n771 VGND.n162 292.5
R3917 VGND.n228 VGND.n225 292.5
R3918 VGND.n262 VGND.n225 292.5
R3919 VGND.n223 VGND.n222 292.5
R3920 VGND.n262 VGND.n223 292.5
R3921 VGND.n858 VGND.n165 288.961
R3922 VGND.n1759 VGND.n141 288.961
R3923 VGND.n258 VGND.n216 288.961
R3924 VGND.n252 VGND.n251 288.961
R3925 VGND.n263 VGND.t200 285.123
R3926 VGND.n1236 VGND.n1235 281.135
R3927 VGND.n1386 VGND.n1385 281.135
R3928 VGND.n1376 VGND.n1375 281.135
R3929 VGND.n1351 VGND.n1350 281.135
R3930 VGND.n1326 VGND.n1325 281.135
R3931 VGND.n1301 VGND.n1300 281.135
R3932 VGND.n1176 VGND.n519 281.135
R3933 VGND.n536 VGND.n529 281.135
R3934 VGND.t368 VGND.t370 275.329
R3935 VGND.n262 VGND.n261 258.13
R3936 VGND.n1001 VGND.n999 257.264
R3937 VGND.n151 VGND.t296 254.272
R3938 VGND.t21 VGND.t23 246.464
R3939 VGND.n565 VGND.t158 230.401
R3940 VGND.n1036 VGND.n1034 226.917
R3941 VGND.n1750 VGND.n165 223.68
R3942 VGND.n1759 VGND.n1758 223.68
R3943 VGND.n258 VGND.n257 223.68
R3944 VGND.n253 VGND.n252 223.68
R3945 VGND.n1763 VGND.n1762 220.702
R3946 VGND.t81 VGND.t363 209.071
R3947 VGND.t363 VGND.t188 209.071
R3948 VGND.t23 VGND.t270 209.071
R3949 VGND.n858 VGND.n163 205.69
R3950 VGND.n156 VGND.n141 205.69
R3951 VGND.n266 VGND.n216 205.69
R3952 VGND.n251 VGND.n232 205.69
R3953 VGND.n1728 VGND.n514 200.744
R3954 VGND.n1303 VGND.n1302 200.744
R3955 VGND.n1328 VGND.n1327 200.744
R3956 VGND.n1353 VGND.n1352 200.744
R3957 VGND.n1378 VGND.n1377 200.744
R3958 VGND.n1387 VGND.n1223 200.744
R3959 VGND.n1260 VGND.n1237 200.744
R3960 VGND.n1724 VGND.n1723 200.744
R3961 VGND.n1028 VGND.n166 196.581
R3962 VGND.n1793 VGND.n1792 195.292
R3963 VGND.n89 VGND.n88 195
R3964 VGND.n88 VGND.n80 195
R3965 VGND.n95 VGND.n94 195
R3966 VGND.n94 VGND.n80 195
R3967 VGND.n101 VGND.n100 195
R3968 VGND.n100 VGND.n80 195
R3969 VGND.n107 VGND.n106 195
R3970 VGND.n106 VGND.n80 195
R3971 VGND.n113 VGND.n112 195
R3972 VGND.n112 VGND.n80 195
R3973 VGND.n119 VGND.n118 195
R3974 VGND.n118 VGND.n80 195
R3975 VGND.n125 VGND.n124 195
R3976 VGND.n124 VGND.n80 195
R3977 VGND.n1774 VGND.n1773 195
R3978 VGND.n1773 VGND.n80 195
R3979 VGND.n86 VGND.n84 195
R3980 VGND.n84 VGND.n80 195
R3981 VGND.n21 VGND.n20 195
R3982 VGND.n20 VGND.n11 195
R3983 VGND.n27 VGND.n26 195
R3984 VGND.n26 VGND.n11 195
R3985 VGND.n33 VGND.n32 195
R3986 VGND.n32 VGND.n11 195
R3987 VGND.n39 VGND.n38 195
R3988 VGND.n38 VGND.n11 195
R3989 VGND.n45 VGND.n44 195
R3990 VGND.n44 VGND.n11 195
R3991 VGND.n51 VGND.n50 195
R3992 VGND.n50 VGND.n11 195
R3993 VGND.n57 VGND.n56 195
R3994 VGND.n56 VGND.n11 195
R3995 VGND.n63 VGND.n62 195
R3996 VGND.n62 VGND.n11 195
R3997 VGND.n1805 VGND.n1804 195
R3998 VGND.n1804 VGND.n11 195
R3999 VGND.n369 VGND.n368 195
R4000 VGND.n368 VGND.n354 195
R4001 VGND.n367 VGND.n366 195
R4002 VGND.n366 VGND.n354 195
R4003 VGND.n377 VGND.n376 195
R4004 VGND.n376 VGND.n354 195
R4005 VGND.n383 VGND.n382 195
R4006 VGND.n382 VGND.n354 195
R4007 VGND.n389 VGND.n388 195
R4008 VGND.n388 VGND.n354 195
R4009 VGND.n395 VGND.n394 195
R4010 VGND.n394 VGND.n354 195
R4011 VGND.n401 VGND.n400 195
R4012 VGND.n400 VGND.n354 195
R4013 VGND.n407 VGND.n406 195
R4014 VGND.n406 VGND.n354 195
R4015 VGND.n413 VGND.n412 195
R4016 VGND.n412 VGND.n354 195
R4017 VGND.n419 VGND.n418 195
R4018 VGND.n418 VGND.n354 195
R4019 VGND.n425 VGND.n424 195
R4020 VGND.n424 VGND.n354 195
R4021 VGND.n431 VGND.n430 195
R4022 VGND.n430 VGND.n354 195
R4023 VGND.n437 VGND.n436 195
R4024 VGND.n436 VGND.n354 195
R4025 VGND.n443 VGND.n442 195
R4026 VGND.n442 VGND.n354 195
R4027 VGND.n449 VGND.n448 195
R4028 VGND.n448 VGND.n354 195
R4029 VGND.n455 VGND.n454 195
R4030 VGND.n454 VGND.n354 195
R4031 VGND.n461 VGND.n460 195
R4032 VGND.n460 VGND.n354 195
R4033 VGND.n467 VGND.n466 195
R4034 VGND.n466 VGND.n354 195
R4035 VGND.n471 VGND.n470 195
R4036 VGND.n470 VGND.n354 195
R4037 VGND.n343 VGND.n340 195
R4038 VGND.n354 VGND.n343 195
R4039 VGND.n872 VGND.n752 195
R4040 VGND.n990 VGND.n752 195
R4041 VGND.n854 VGND.n753 195
R4042 VGND.n990 VGND.n753 195
R4043 VGND.n877 VGND.n751 195
R4044 VGND.n990 VGND.n751 195
R4045 VGND.n851 VGND.n754 195
R4046 VGND.n990 VGND.n754 195
R4047 VGND.n894 VGND.n750 195
R4048 VGND.n990 VGND.n750 195
R4049 VGND.n840 VGND.n755 195
R4050 VGND.n990 VGND.n755 195
R4051 VGND.n899 VGND.n749 195
R4052 VGND.n990 VGND.n749 195
R4053 VGND.n837 VGND.n756 195
R4054 VGND.n990 VGND.n756 195
R4055 VGND.n916 VGND.n748 195
R4056 VGND.n990 VGND.n748 195
R4057 VGND.n826 VGND.n757 195
R4058 VGND.n990 VGND.n757 195
R4059 VGND.n921 VGND.n747 195
R4060 VGND.n990 VGND.n747 195
R4061 VGND.n823 VGND.n758 195
R4062 VGND.n990 VGND.n758 195
R4063 VGND.n938 VGND.n746 195
R4064 VGND.n990 VGND.n746 195
R4065 VGND.n812 VGND.n759 195
R4066 VGND.n990 VGND.n759 195
R4067 VGND.n943 VGND.n745 195
R4068 VGND.n990 VGND.n745 195
R4069 VGND.n809 VGND.n760 195
R4070 VGND.n990 VGND.n760 195
R4071 VGND.n960 VGND.n744 195
R4072 VGND.n990 VGND.n744 195
R4073 VGND.n798 VGND.n761 195
R4074 VGND.n990 VGND.n761 195
R4075 VGND.n965 VGND.n743 195
R4076 VGND.n990 VGND.n743 195
R4077 VGND.n795 VGND.n762 195
R4078 VGND.n990 VGND.n762 195
R4079 VGND.n765 VGND.n742 195
R4080 VGND.n990 VGND.n742 195
R4081 VGND.n988 VGND.n987 195
R4082 VGND.n990 VGND.n988 195
R4083 VGND.n992 VGND.n991 195
R4084 VGND.n991 VGND.n990 195
R4085 VGND.n989 VGND.n738 195
R4086 VGND.n990 VGND.n989 195
R4087 VGND.n150 VGND.n149 195
R4088 VGND.n151 VGND.n150 195
R4089 VGND.n153 VGND.n152 195
R4090 VGND.n152 VGND.n151 195
R4091 VGND.n243 VGND.n242 195
R4092 VGND.n242 VGND.n241 195
R4093 VGND.n240 VGND.n235 195
R4094 VGND.n241 VGND.n240 195
R4095 VGND.n272 VGND.n207 195
R4096 VGND.n301 VGND.n207 195
R4097 VGND.n213 VGND.n209 195
R4098 VGND.n301 VGND.n209 195
R4099 VGND.n212 VGND.n206 195
R4100 VGND.n301 VGND.n206 195
R4101 VGND.n281 VGND.n280 195
R4102 VGND.n301 VGND.n281 195
R4103 VGND.n291 VGND.n205 195
R4104 VGND.n301 VGND.n205 195
R4105 VGND.n286 VGND.n282 195
R4106 VGND.n301 VGND.n282 195
R4107 VGND.n285 VGND.n204 195
R4108 VGND.n301 VGND.n204 195
R4109 VGND.n300 VGND.n299 195
R4110 VGND.n301 VGND.n300 195
R4111 VGND.t370 VGND.t372 191.115
R4112 VGND.n186 VGND.n184 190.601
R4113 VGND.n1209 VGND.n1208 184.73
R4114 VGND.n1299 VGND.n1285 184.73
R4115 VGND.n1324 VGND.n1310 184.73
R4116 VGND.n1349 VGND.n1335 184.73
R4117 VGND.n1374 VGND.n1360 184.73
R4118 VGND.n1390 VGND.n1389 184.73
R4119 VGND.n1247 VGND.n1246 184.73
R4120 VGND.n1722 VGND.n533 184.73
R4121 VGND VGND.n728 161.595
R4122 VGND VGND.n171 161.595
R4123 VGND.n1726 VGND.n524 155.677
R4124 VGND.n1728 VGND.n517 152.744
R4125 VGND.n1303 VGND.n1277 152.744
R4126 VGND.n1328 VGND.n1274 152.744
R4127 VGND.n1353 VGND.n1271 152.744
R4128 VGND.n1378 VGND.n1268 152.744
R4129 VGND.n1234 VGND.n1223 152.744
R4130 VGND.n1260 VGND.n1259 152.744
R4131 VGND.n1724 VGND.n530 152.744
R4132 VGND.t372 VGND.n1794 149.852
R4133 VGND.n509 VGND.n354 146.72
R4134 VGND.n1534 VGND.n1523 146.25
R4135 VGND.n1535 VGND.n1534 146.25
R4136 VGND.n1545 VGND.n1544 146.25
R4137 VGND.n1546 VGND.n1545 146.25
R4138 VGND.n1411 VGND.n1410 146.25
R4139 VGND.n1410 VGND.n1409 146.25
R4140 VGND.n1419 VGND.n1412 146.25
R4141 VGND.n1420 VGND.n1419 146.25
R4142 VGND.n1511 VGND.n1423 146.25
R4143 VGND.n1423 VGND.n1422 146.25
R4144 VGND.n1431 VGND.n1424 146.25
R4145 VGND.n1432 VGND.n1431 146.25
R4146 VGND.n1502 VGND.n1435 146.25
R4147 VGND.n1435 VGND.n1434 146.25
R4148 VGND.n1443 VGND.n1436 146.25
R4149 VGND.n1444 VGND.n1443 146.25
R4150 VGND.n1493 VGND.n1447 146.25
R4151 VGND.n1447 VGND.n1446 146.25
R4152 VGND.n1455 VGND.n1448 146.25
R4153 VGND.n1456 VGND.n1455 146.25
R4154 VGND.n1484 VGND.n1459 146.25
R4155 VGND.n1459 VGND.n1458 146.25
R4156 VGND.n1467 VGND.n1460 146.25
R4157 VGND.n1468 VGND.n1467 146.25
R4158 VGND.n1475 VGND.n1471 146.25
R4159 VGND.n1471 VGND.n1470 146.25
R4160 VGND.n1552 VGND.n1551 146.25
R4161 VGND.n1551 VGND.n1550 146.25
R4162 VGND.n1160 VGND.n1150 146.25
R4163 VGND.n1161 VGND.n1160 146.25
R4164 VGND.n1149 VGND.n1148 146.25
R4165 VGND.n1148 VGND.n1147 146.25
R4166 VGND.n1566 VGND.n1565 146.25
R4167 VGND.n1567 VGND.n1566 146.25
R4168 VGND.n1707 VGND.n1706 146.25
R4169 VGND.n1708 VGND.n1707 146.25
R4170 VGND.n1532 VGND.n1531 146.25
R4171 VGND.n1532 VGND.n555 146.25
R4172 VGND.n1654 VGND.n74 146.25
R4173 VGND.n1655 VGND.n1654 146.25
R4174 VGND.n1658 VGND.n1657 146.25
R4175 VGND.n1657 VGND.n1656 146.25
R4176 VGND.n1651 VGND.n1634 146.25
R4177 VGND.n1652 VGND.n1651 146.25
R4178 VGND.n1649 VGND.n1633 146.25
R4179 VGND.n1650 VGND.n1649 146.25
R4180 VGND.n1672 VGND.n1671 146.25
R4181 VGND.n1673 VGND.n1672 146.25
R4182 VGND.n1676 VGND.n1675 146.25
R4183 VGND.n1675 VGND.n1674 146.25
R4184 VGND.n1624 VGND.n1610 146.25
R4185 VGND.n1625 VGND.n1624 146.25
R4186 VGND.n1622 VGND.n1609 146.25
R4187 VGND.n1623 VGND.n1622 146.25
R4188 VGND.n1690 VGND.n1689 146.25
R4189 VGND.n1691 VGND.n1690 146.25
R4190 VGND.n1694 VGND.n1693 146.25
R4191 VGND.n1693 VGND.n1692 146.25
R4192 VGND.n1600 VGND.n1586 146.25
R4193 VGND.n1601 VGND.n1600 146.25
R4194 VGND.n1598 VGND.n1585 146.25
R4195 VGND.n1599 VGND.n1598 146.25
R4196 VGND.n1792 VGND.n69 146.25
R4197 VGND.n1775 VGND.n79 146.25
R4198 VGND.n1791 VGND.n79 146.25
R4199 VGND.n1777 VGND.n81 146.25
R4200 VGND.n1791 VGND.n81 146.25
R4201 VGND.n1779 VGND.n78 146.25
R4202 VGND.n1791 VGND.n78 146.25
R4203 VGND.n1781 VGND.n82 146.25
R4204 VGND.n1791 VGND.n82 146.25
R4205 VGND.n1783 VGND.n77 146.25
R4206 VGND.n1791 VGND.n77 146.25
R4207 VGND.n1785 VGND.n83 146.25
R4208 VGND.n1791 VGND.n83 146.25
R4209 VGND.n1787 VGND.n76 146.25
R4210 VGND.n1791 VGND.n76 146.25
R4211 VGND.n1790 VGND.n1789 146.25
R4212 VGND.n1791 VGND.n1790 146.25
R4213 VGND.n1806 VGND.n12 146.25
R4214 VGND.n1824 VGND.n12 146.25
R4215 VGND.n1808 VGND.n10 146.25
R4216 VGND.n1824 VGND.n10 146.25
R4217 VGND.n1810 VGND.n13 146.25
R4218 VGND.n1824 VGND.n13 146.25
R4219 VGND.n1812 VGND.n9 146.25
R4220 VGND.n1824 VGND.n9 146.25
R4221 VGND.n1814 VGND.n14 146.25
R4222 VGND.n1824 VGND.n14 146.25
R4223 VGND.n1816 VGND.n8 146.25
R4224 VGND.n1824 VGND.n8 146.25
R4225 VGND.n1818 VGND.n15 146.25
R4226 VGND.n1824 VGND.n15 146.25
R4227 VGND.n1820 VGND.n7 146.25
R4228 VGND.n1824 VGND.n7 146.25
R4229 VGND.n1823 VGND.n1822 146.25
R4230 VGND.n1824 VGND.n1823 146.25
R4231 VGND.n475 VGND.n355 146.25
R4232 VGND.n509 VGND.n355 146.25
R4233 VGND.n477 VGND.n353 146.25
R4234 VGND.n509 VGND.n353 146.25
R4235 VGND.n479 VGND.n356 146.25
R4236 VGND.n509 VGND.n356 146.25
R4237 VGND.n481 VGND.n352 146.25
R4238 VGND.n509 VGND.n352 146.25
R4239 VGND.n483 VGND.n357 146.25
R4240 VGND.n509 VGND.n357 146.25
R4241 VGND.n485 VGND.n351 146.25
R4242 VGND.n509 VGND.n351 146.25
R4243 VGND.n487 VGND.n358 146.25
R4244 VGND.n509 VGND.n358 146.25
R4245 VGND.n489 VGND.n350 146.25
R4246 VGND.n509 VGND.n350 146.25
R4247 VGND.n491 VGND.n359 146.25
R4248 VGND.n509 VGND.n359 146.25
R4249 VGND.n493 VGND.n349 146.25
R4250 VGND.n509 VGND.n349 146.25
R4251 VGND.n495 VGND.n360 146.25
R4252 VGND.n509 VGND.n360 146.25
R4253 VGND.n497 VGND.n348 146.25
R4254 VGND.n509 VGND.n348 146.25
R4255 VGND.n499 VGND.n361 146.25
R4256 VGND.n509 VGND.n361 146.25
R4257 VGND.n501 VGND.n347 146.25
R4258 VGND.n509 VGND.n347 146.25
R4259 VGND.n503 VGND.n362 146.25
R4260 VGND.n509 VGND.n362 146.25
R4261 VGND.n505 VGND.n346 146.25
R4262 VGND.n509 VGND.n346 146.25
R4263 VGND.n508 VGND.n507 146.25
R4264 VGND.n509 VGND.n508 146.25
R4265 VGND.n371 VGND.n345 146.25
R4266 VGND.n509 VGND.n345 146.25
R4267 VGND.n511 VGND.n510 146.25
R4268 VGND.n510 VGND.n509 146.25
R4269 VGND.n1756 VGND.n1755 146.25
R4270 VGND.n1755 VGND.n1754 146.25
R4271 VGND.n1753 VGND.n1752 146.25
R4272 VGND.n1754 VGND.n1753 146.25
R4273 VGND.n873 VGND.n856 146.25
R4274 VGND.n856 VGND.n771 146.25
R4275 VGND.n878 VGND.n853 146.25
R4276 VGND.n853 VGND.n771 146.25
R4277 VGND.n882 VGND.n780 146.25
R4278 VGND.n976 VGND.n780 146.25
R4279 VGND.n846 VGND.n782 146.25
R4280 VGND.n976 VGND.n782 146.25
R4281 VGND.n888 VGND.n779 146.25
R4282 VGND.n976 VGND.n779 146.25
R4283 VGND.n843 VGND.n783 146.25
R4284 VGND.n976 VGND.n783 146.25
R4285 VGND.n895 VGND.n842 146.25
R4286 VGND.n842 VGND.n771 146.25
R4287 VGND.n900 VGND.n839 146.25
R4288 VGND.n839 VGND.n771 146.25
R4289 VGND.n904 VGND.n778 146.25
R4290 VGND.n976 VGND.n778 146.25
R4291 VGND.n832 VGND.n784 146.25
R4292 VGND.n976 VGND.n784 146.25
R4293 VGND.n910 VGND.n777 146.25
R4294 VGND.n976 VGND.n777 146.25
R4295 VGND.n829 VGND.n785 146.25
R4296 VGND.n976 VGND.n785 146.25
R4297 VGND.n917 VGND.n828 146.25
R4298 VGND.n828 VGND.n771 146.25
R4299 VGND.n922 VGND.n825 146.25
R4300 VGND.n825 VGND.n771 146.25
R4301 VGND.n926 VGND.n776 146.25
R4302 VGND.n976 VGND.n776 146.25
R4303 VGND.n818 VGND.n786 146.25
R4304 VGND.n976 VGND.n786 146.25
R4305 VGND.n932 VGND.n775 146.25
R4306 VGND.n976 VGND.n775 146.25
R4307 VGND.n815 VGND.n787 146.25
R4308 VGND.n976 VGND.n787 146.25
R4309 VGND.n939 VGND.n814 146.25
R4310 VGND.n814 VGND.n771 146.25
R4311 VGND.n944 VGND.n811 146.25
R4312 VGND.n811 VGND.n771 146.25
R4313 VGND.n948 VGND.n774 146.25
R4314 VGND.n976 VGND.n774 146.25
R4315 VGND.n804 VGND.n788 146.25
R4316 VGND.n976 VGND.n788 146.25
R4317 VGND.n954 VGND.n773 146.25
R4318 VGND.n976 VGND.n773 146.25
R4319 VGND.n801 VGND.n789 146.25
R4320 VGND.n976 VGND.n789 146.25
R4321 VGND.n961 VGND.n800 146.25
R4322 VGND.n800 VGND.n771 146.25
R4323 VGND.n966 VGND.n797 146.25
R4324 VGND.n797 VGND.n771 146.25
R4325 VGND.n794 VGND.n772 146.25
R4326 VGND.n976 VGND.n772 146.25
R4327 VGND.n974 VGND.n973 146.25
R4328 VGND.n976 VGND.n974 146.25
R4329 VGND.n978 VGND.n977 146.25
R4330 VGND.n977 VGND.n976 146.25
R4331 VGND.n975 VGND.n766 146.25
R4332 VGND.n976 VGND.n975 146.25
R4333 VGND.n764 VGND.n763 146.25
R4334 VGND.n771 VGND.n763 146.25
R4335 VGND.n993 VGND.n740 146.25
R4336 VGND.n771 VGND.n740 146.25
R4337 VGND.n1007 VGND.n1006 146.25
R4338 VGND.n1006 VGND.n1005 146.25
R4339 VGND.n1000 VGND.n733 146.25
R4340 VGND.n1001 VGND.n1000 146.25
R4341 VGND.n998 VGND.n732 146.25
R4342 VGND.n999 VGND.n998 146.25
R4343 VGND.n1016 VGND.n1015 146.25
R4344 VGND.n1017 VGND.n1016 146.25
R4345 VGND.n145 VGND.n144 146.25
R4346 VGND.n146 VGND.n145 146.25
R4347 VGND.n244 VGND.n237 146.25
R4348 VGND.n238 VGND.n237 146.25
R4349 VGND.n231 VGND.n224 146.25
R4350 VGND.n263 VGND.n224 146.25
R4351 VGND.n265 VGND.n264 146.25
R4352 VGND.n264 VGND.n263 146.25
R4353 VGND.n273 VGND.n215 146.25
R4354 VGND.n215 VGND.n191 146.25
R4355 VGND.n211 VGND.n210 146.25
R4356 VGND.n210 VGND.n191 146.25
R4357 VGND.n305 VGND.n304 146.25
R4358 VGND.n304 VGND.n303 146.25
R4359 VGND.n302 VGND.n199 146.25
R4360 VGND.n303 VGND.n302 146.25
R4361 VGND.n195 VGND.n193 146.25
R4362 VGND.n303 VGND.n193 146.25
R4363 VGND.n194 VGND.n192 146.25
R4364 VGND.n303 VGND.n192 146.25
R4365 VGND.n292 VGND.n288 146.25
R4366 VGND.n288 VGND.n191 146.25
R4367 VGND.n284 VGND.n283 146.25
R4368 VGND.n283 VGND.n191 146.25
R4369 VGND.n319 VGND.n318 146.25
R4370 VGND.n318 VGND.n317 146.25
R4371 VGND.n185 VGND.n176 146.25
R4372 VGND.n186 VGND.n185 146.25
R4373 VGND.n183 VGND.n175 146.25
R4374 VGND.n184 VGND.n183 146.25
R4375 VGND.n328 VGND.n327 146.25
R4376 VGND.n329 VGND.n328 146.25
R4377 VGND.n1751 VGND.n1750 143.361
R4378 VGND.n1758 VGND.n142 143.361
R4379 VGND.n257 VGND.n222 143.361
R4380 VGND.n253 VGND.n228 143.361
R4381 VGND.n606 VGND.n592 141.846
R4382 VGND.n630 VGND.n616 141.846
R4383 VGND.n654 VGND.n640 141.846
R4384 VGND.n678 VGND.n664 141.846
R4385 VGND.n696 VGND.n688 141.846
R4386 VGND.n315 VGND.n314 141.596
R4387 VGND.n608 VGND.n606 141.343
R4388 VGND.n632 VGND.n630 141.343
R4389 VGND.n656 VGND.n654 141.343
R4390 VGND.n680 VGND.n678 141.343
R4391 VGND.n698 VGND.n696 141.343
R4392 VGND.n1005 VGND.n1004 140.327
R4393 VGND.t74 VGND.n208 135.933
R4394 VGND.n1020 VGND.n1018 135.099
R4395 VGND.n1797 VGND.n69 133.755
R4396 VGND.n1797 VGND.n74 133.755
R4397 VGND.n1659 VGND.n1658 133.755
R4398 VGND.n1659 VGND.n1634 133.755
R4399 VGND.n1633 VGND.n1628 133.755
R4400 VGND.n1671 VGND.n1628 133.755
R4401 VGND.n1677 VGND.n1676 133.755
R4402 VGND.n1677 VGND.n1610 133.755
R4403 VGND.n1609 VGND.n1604 133.755
R4404 VGND.n1689 VGND.n1604 133.755
R4405 VGND.n1695 VGND.n1694 133.755
R4406 VGND.n1695 VGND.n1586 133.755
R4407 VGND.n1585 VGND.n1580 133.755
R4408 VGND.n1706 VGND.n1580 133.755
R4409 VGND.n1538 VGND.n1531 133.755
R4410 VGND.n1538 VGND.n1523 133.755
R4411 VGND.n1544 VGND.n1402 133.755
R4412 VGND.n1411 VGND.n1402 133.755
R4413 VGND.n1512 VGND.n1412 133.755
R4414 VGND.n1512 VGND.n1511 133.755
R4415 VGND.n1503 VGND.n1424 133.755
R4416 VGND.n1503 VGND.n1502 133.755
R4417 VGND.n1494 VGND.n1436 133.755
R4418 VGND.n1494 VGND.n1493 133.755
R4419 VGND.n1485 VGND.n1448 133.755
R4420 VGND.n1485 VGND.n1484 133.755
R4421 VGND.n1476 VGND.n1460 133.755
R4422 VGND.n1476 VGND.n1475 133.755
R4423 VGND.n1553 VGND.n1552 133.755
R4424 VGND.n1553 VGND.n1150 133.755
R4425 VGND.n1149 VGND.n567 133.755
R4426 VGND.n1565 VGND.n567 133.755
R4427 VGND.n241 VGND.n239 133.377
R4428 VGND.n1211 VGND.n1210 131.84
R4429 VGND.n1287 VGND.n1286 131.84
R4430 VGND.n1312 VGND.n1311 131.84
R4431 VGND.n1337 VGND.n1336 131.84
R4432 VGND.n1362 VGND.n1361 131.84
R4433 VGND.n1392 VGND.n1391 131.84
R4434 VGND.n1248 VGND.n1242 131.84
R4435 VGND.n1397 VGND.n1396 131.84
R4436 VGND.n1206 VGND.n1205 125.35
R4437 VGND.n1289 VGND.n1288 125.35
R4438 VGND.n1314 VGND.n1313 125.35
R4439 VGND.n1339 VGND.n1338 125.35
R4440 VGND.n1364 VGND.n1363 125.35
R4441 VGND.n1229 VGND.n1222 125.35
R4442 VGND.n1250 VGND.n1249 125.35
R4443 VGND.n1398 VGND.n554 125.35
R4444 VGND.n255 VGND.t30 123.16
R4445 VGND.n313 VGND.n191 118.132
R4446 VGND.n1715 VGND.n1714 117.001
R4447 VGND.n1714 VGND.n1713 117.001
R4448 VGND.n1202 VGND.n1201 117.001
R4449 VGND.n1202 VGND.n545 117.001
R4450 VGND.n1207 VGND.n544 117.001
R4451 VGND.n1719 VGND.n544 117.001
R4452 VGND.n1294 VGND.n1293 117.001
R4453 VGND.n1293 VGND.n545 117.001
R4454 VGND.n1298 VGND.n543 117.001
R4455 VGND.n1719 VGND.n543 117.001
R4456 VGND.n1319 VGND.n1318 117.001
R4457 VGND.n1318 VGND.n545 117.001
R4458 VGND.n1323 VGND.n542 117.001
R4459 VGND.n1719 VGND.n542 117.001
R4460 VGND.n1344 VGND.n1343 117.001
R4461 VGND.n1343 VGND.n545 117.001
R4462 VGND.n1348 VGND.n541 117.001
R4463 VGND.n1719 VGND.n541 117.001
R4464 VGND.n1369 VGND.n1368 117.001
R4465 VGND.n1368 VGND.n545 117.001
R4466 VGND.n1373 VGND.n540 117.001
R4467 VGND.n1719 VGND.n540 117.001
R4468 VGND.n1233 VGND.n1232 117.001
R4469 VGND.n1232 VGND.n545 117.001
R4470 VGND.n1388 VGND.n539 117.001
R4471 VGND.n1719 VGND.n539 117.001
R4472 VGND.n1254 VGND.n1253 117.001
R4473 VGND.n1253 VGND.n545 117.001
R4474 VGND.n1245 VGND.n538 117.001
R4475 VGND.n1719 VGND.n538 117.001
R4476 VGND.n1721 VGND.n1720 117.001
R4477 VGND.n1720 VGND.n1719 117.001
R4478 VGND.t437 VGND.t546 115.859
R4479 VGND.n1824 VGND.n11 114.246
R4480 VGND.n1017 VGND.t474 112.261
R4481 VGND.n999 VGND.t18 112.261
R4482 VGND.t482 VGND.n1001 112.261
R4483 VGND.n1005 VGND.t399 112.261
R4484 VGND.n1211 VGND.n1198 111.68
R4485 VGND.n1297 VGND.n1286 111.68
R4486 VGND.n1322 VGND.n1311 111.68
R4487 VGND.n1347 VGND.n1336 111.68
R4488 VGND.n1372 VGND.n1361 111.68
R4489 VGND.n1392 VGND.n1221 111.68
R4490 VGND.n1244 VGND.n1242 111.68
R4491 VGND.n1396 VGND.n534 111.68
R4492 VGND.n1710 VGND.n1709 111.663
R4493 VGND.n1833 VGND.n1 110.933
R4494 VGND.n1833 VGND.n1832 110.933
R4495 VGND.n1765 VGND.n130 110.933
R4496 VGND.n1765 VGND.n132 110.933
R4497 VGND.n320 VGND.n176 105.695
R4498 VGND.n320 VGND.n319 105.695
R4499 VGND.n311 VGND.n194 105.695
R4500 VGND.n311 VGND.n195 105.695
R4501 VGND.n306 VGND.n199 105.695
R4502 VGND.n306 VGND.n305 105.695
R4503 VGND.n1008 VGND.n733 105.695
R4504 VGND.n1008 VGND.n1007 105.695
R4505 VGND.n979 VGND.n766 105.695
R4506 VGND.n979 VGND.n978 105.695
R4507 VGND.n973 VGND.n791 105.695
R4508 VGND.n794 VGND.n791 105.695
R4509 VGND.n955 VGND.n801 105.695
R4510 VGND.n955 VGND.n954 105.695
R4511 VGND.n949 VGND.n804 105.695
R4512 VGND.n949 VGND.n948 105.695
R4513 VGND.n933 VGND.n815 105.695
R4514 VGND.n933 VGND.n932 105.695
R4515 VGND.n927 VGND.n818 105.695
R4516 VGND.n927 VGND.n926 105.695
R4517 VGND.n911 VGND.n829 105.695
R4518 VGND.n911 VGND.n910 105.695
R4519 VGND.n905 VGND.n832 105.695
R4520 VGND.n905 VGND.n904 105.695
R4521 VGND.n889 VGND.n843 105.695
R4522 VGND.n889 VGND.n888 105.695
R4523 VGND.n883 VGND.n846 105.695
R4524 VGND.n883 VGND.n882 105.695
R4525 VGND.n732 VGND.n727 105.695
R4526 VGND.n1015 VGND.n727 105.695
R4527 VGND.n175 VGND.n170 105.695
R4528 VGND.n327 VGND.n170 105.695
R4529 VGND.n317 VGND.n316 103.965
R4530 VGND.n1794 VGND.t28 102.638
R4531 VGND.n1201 VGND.n517 101.555
R4532 VGND.n1294 VGND.n1277 101.555
R4533 VGND.n1319 VGND.n1274 101.555
R4534 VGND.n1344 VGND.n1271 101.555
R4535 VGND.n1369 VGND.n1268 101.555
R4536 VGND.n1234 VGND.n1233 101.555
R4537 VGND.n1259 VGND.n1254 101.555
R4538 VGND.n1715 VGND.n530 101.555
R4539 VGND.n1004 VGND.n1003 99.0083
R4540 VGND.n1199 VGND.n546 97.5005
R4541 VGND.n1719 VGND.n546 97.5005
R4542 VGND.n1206 VGND.n1178 97.5005
R4543 VGND.n1400 VGND.n1178 97.5005
R4544 VGND.n1209 VGND.n1177 97.5005
R4545 VGND.n1400 VGND.n1177 97.5005
R4546 VGND.n1296 VGND.n547 97.5005
R4547 VGND.n1719 VGND.n547 97.5005
R4548 VGND.n1288 VGND.n1179 97.5005
R4549 VGND.n1400 VGND.n1179 97.5005
R4550 VGND.n1285 VGND.n1175 97.5005
R4551 VGND.n1400 VGND.n1175 97.5005
R4552 VGND.n1321 VGND.n548 97.5005
R4553 VGND.n1719 VGND.n548 97.5005
R4554 VGND.n1313 VGND.n1180 97.5005
R4555 VGND.n1400 VGND.n1180 97.5005
R4556 VGND.n1310 VGND.n1174 97.5005
R4557 VGND.n1400 VGND.n1174 97.5005
R4558 VGND.n1346 VGND.n549 97.5005
R4559 VGND.n1719 VGND.n549 97.5005
R4560 VGND.n1338 VGND.n1181 97.5005
R4561 VGND.n1400 VGND.n1181 97.5005
R4562 VGND.n1335 VGND.n1173 97.5005
R4563 VGND.n1400 VGND.n1173 97.5005
R4564 VGND.n1371 VGND.n550 97.5005
R4565 VGND.n1719 VGND.n550 97.5005
R4566 VGND.n1363 VGND.n1182 97.5005
R4567 VGND.n1400 VGND.n1182 97.5005
R4568 VGND.n1360 VGND.n1172 97.5005
R4569 VGND.n1400 VGND.n1172 97.5005
R4570 VGND.n1227 VGND.n551 97.5005
R4571 VGND.n1719 VGND.n551 97.5005
R4572 VGND.n1222 VGND.n1183 97.5005
R4573 VGND.n1400 VGND.n1183 97.5005
R4574 VGND.n1390 VGND.n1171 97.5005
R4575 VGND.n1400 VGND.n1171 97.5005
R4576 VGND.n1243 VGND.n552 97.5005
R4577 VGND.n1719 VGND.n552 97.5005
R4578 VGND.n1249 VGND.n1184 97.5005
R4579 VGND.n1400 VGND.n1184 97.5005
R4580 VGND.n1247 VGND.n1170 97.5005
R4581 VGND.n1400 VGND.n1170 97.5005
R4582 VGND.n1718 VGND.n1717 97.5005
R4583 VGND.n1719 VGND.n1718 97.5005
R4584 VGND.n1399 VGND.n1398 97.5005
R4585 VGND.n1400 VGND.n1399 97.5005
R4586 VGND.n1169 VGND.n533 97.5005
R4587 VGND.n1400 VGND.n1169 97.5005
R4588 VGND.n134 VGND.n130 97.5005
R4589 VGND.n1762 VGND.n134 97.5005
R4590 VGND.n133 VGND.n132 97.5005
R4591 VGND.n1762 VGND.n133 97.5005
R4592 VGND.n1832 VGND.n1831 97.5005
R4593 VGND.n1831 VGND.n1830 97.5005
R4594 VGND.n1829 VGND.n1 97.5005
R4595 VGND.n1830 VGND.n1829 97.5005
R4596 VGND.n1752 VGND.n1751 93.4405
R4597 VGND.n1756 VGND.n142 93.4405
R4598 VGND.n265 VGND.n222 93.4405
R4599 VGND.n231 VGND.n228 93.4405
R4600 VGND.n1794 VGND.n1793 93.0698
R4601 VGND.n1400 VGND.n1168 90.9633
R4602 VGND.n1825 VGND.n6 87.9761
R4603 VGND.n1735 VGND.t349 84.5161
R4604 VGND.n1045 VGND.t342 84.5161
R4605 VGND.n1030 VGND.t195 84.5161
R4606 VGND.n1058 VGND.t238 84.5161
R4607 VGND.n1063 VGND.t129 84.5161
R4608 VGND.n701 VGND.t96 84.5161
R4609 VGND.n690 VGND.t14 84.5161
R4610 VGND.n1084 VGND.t340 84.5161
R4611 VGND.n666 VGND.t533 84.5161
R4612 VGND.n1097 VGND.t484 84.5161
R4613 VGND.n642 VGND.t8 84.5161
R4614 VGND.n1110 VGND.t257 84.5161
R4615 VGND.n618 VGND.t471 84.5161
R4616 VGND.n1123 VGND.t460 84.5161
R4617 VGND.n594 VGND.t36 84.5161
R4618 VGND.n1136 VGND.t202 84.5161
R4619 VGND.n236 VGND.t295 84.1574
R4620 VGND.n214 VGND.t402 84.1574
R4621 VGND.n277 VGND.t426 84.1574
R4622 VGND.n287 VGND.t409 84.1574
R4623 VGND.n296 VGND.t75 84.1574
R4624 VGND.n147 VGND.t297 84.1574
R4625 VGND.n855 VGND.t187 84.1574
R4626 VGND.n852 VGND.t548 84.1574
R4627 VGND.n841 VGND.t125 84.1574
R4628 VGND.n838 VGND.t560 84.1574
R4629 VGND.n827 VGND.t534 84.1574
R4630 VGND.n824 VGND.t130 84.1574
R4631 VGND.n813 VGND.t524 84.1574
R4632 VGND.n810 VGND.t481 84.1574
R4633 VGND.n799 VGND.t223 84.1574
R4634 VGND.n796 VGND.t241 84.1574
R4635 VGND.n984 VGND.t410 84.1574
R4636 VGND.n739 VGND.t192 84.1574
R4637 VGND.n129 VGND.t413 84.1574
R4638 VGND.n126 VGND.t149 84.1574
R4639 VGND.n120 VGND.t147 84.1574
R4640 VGND.n114 VGND.t150 84.1574
R4641 VGND.n108 VGND.t148 84.1574
R4642 VGND.n102 VGND.t376 84.1574
R4643 VGND.n96 VGND.t382 84.1574
R4644 VGND.n90 VGND.t379 84.1574
R4645 VGND.n67 VGND.t127 84.1574
R4646 VGND.n64 VGND.t86 84.1574
R4647 VGND.n58 VGND.t554 84.1574
R4648 VGND.n52 VGND.t244 84.1574
R4649 VGND.n46 VGND.t549 84.1574
R4650 VGND.n40 VGND.t94 84.1574
R4651 VGND.n34 VGND.t425 84.1574
R4652 VGND.n28 VGND.t29 84.1574
R4653 VGND.n22 VGND.t526 84.1574
R4654 VGND.n473 VGND.t528 84.1574
R4655 VGND.n468 VGND.t527 84.1574
R4656 VGND.n462 VGND.t525 84.1574
R4657 VGND.n456 VGND.t132 84.1574
R4658 VGND.n450 VGND.t136 84.1574
R4659 VGND.n444 VGND.t280 84.1574
R4660 VGND.n438 VGND.t355 84.1574
R4661 VGND.n432 VGND.t134 84.1574
R4662 VGND.n426 VGND.t133 84.1574
R4663 VGND.n420 VGND.t135 84.1574
R4664 VGND.n414 VGND.t106 84.1574
R4665 VGND.n408 VGND.t137 84.1574
R4666 VGND.n402 VGND.t561 84.1574
R4667 VGND.n396 VGND.t356 84.1574
R4668 VGND.n390 VGND.t163 84.1574
R4669 VGND.n384 VGND.t354 84.1574
R4670 VGND.n378 VGND.t131 84.1574
R4671 VGND.n373 VGND.t180 84.1574
R4672 VGND.n341 VGND.t556 84.1574
R4673 VGND.n201 VGND.t393 83.7172
R4674 VGND.n197 VGND.t320 83.7172
R4675 VGND.n178 VGND.t395 83.7172
R4676 VGND.n174 VGND.t505 83.7172
R4677 VGND.n848 VGND.t362 83.7172
R4678 VGND.n845 VGND.t284 83.7172
R4679 VGND.n834 VGND.t123 83.7172
R4680 VGND.n831 VGND.t358 83.7172
R4681 VGND.n820 VGND.t298 83.7172
R4682 VGND.n817 VGND.t224 83.7172
R4683 VGND.n806 VGND.t261 83.7172
R4684 VGND.n803 VGND.t478 83.7172
R4685 VGND.n793 VGND.t222 83.7172
R4686 VGND.n768 VGND.t204 83.7172
R4687 VGND.n735 VGND.t400 83.7172
R4688 VGND.n731 VGND.t475 83.7172
R4689 VGND.n716 VGND.n704 83.5719
R4690 VGND.n716 VGND.n715 83.5719
R4691 VGND.n718 VGND.n702 83.5719
R4692 VGND.n719 VGND.n718 83.5719
R4693 VGND.n1072 VGND.n1071 83.5719
R4694 VGND.n1071 VGND.n1070 83.5719
R4695 VGND.n1076 VGND.n1075 83.5719
R4696 VGND.n1077 VGND.n1076 83.5719
R4697 VGND.n685 VGND.n672 83.5719
R4698 VGND.n686 VGND.n685 83.5719
R4699 VGND.n676 VGND.n668 83.5719
R4700 VGND.n679 VGND.n676 83.5719
R4701 VGND.n1089 VGND.n1088 83.5719
R4702 VGND.n1090 VGND.n1089 83.5719
R4703 VGND.n661 VGND.n648 83.5719
R4704 VGND.n662 VGND.n661 83.5719
R4705 VGND.n652 VGND.n644 83.5719
R4706 VGND.n655 VGND.n652 83.5719
R4707 VGND.n1102 VGND.n1101 83.5719
R4708 VGND.n1103 VGND.n1102 83.5719
R4709 VGND.n637 VGND.n624 83.5719
R4710 VGND.n638 VGND.n637 83.5719
R4711 VGND.n628 VGND.n620 83.5719
R4712 VGND.n631 VGND.n628 83.5719
R4713 VGND.n1115 VGND.n1114 83.5719
R4714 VGND.n1116 VGND.n1115 83.5719
R4715 VGND.n613 VGND.n600 83.5719
R4716 VGND.n614 VGND.n613 83.5719
R4717 VGND.n604 VGND.n596 83.5719
R4718 VGND.n607 VGND.n604 83.5719
R4719 VGND.n1128 VGND.n1127 83.5719
R4720 VGND.n1129 VGND.n1128 83.5719
R4721 VGND.n589 VGND.n578 83.5719
R4722 VGND.n590 VGND.n589 83.5719
R4723 VGND.n583 VGND.n574 83.5719
R4724 VGND.n583 VGND.n582 83.5719
R4725 VGND.n335 VGND.n334 83.5719
R4726 VGND.n334 VGND.n332 83.5719
R4727 VGND.n1738 VGND.n1737 83.5719
R4728 VGND.n1739 VGND.n1738 83.5719
R4729 VGND.n1043 VGND.n1042 83.5719
R4730 VGND.n1042 VGND.n1041 83.5719
R4731 VGND.n1050 VGND.n1049 83.5719
R4732 VGND.n1051 VGND.n1050 83.5719
R4733 VGND.n1025 VGND.n709 83.5719
R4734 VGND.n1026 VGND.n1025 83.5719
R4735 VGND.n713 VGND.n705 83.5719
R4736 VGND.n1019 VGND.n713 83.5719
R4737 VGND.n184 VGND.t16 83.1719
R4738 VGND.t126 VGND.n186 83.1719
R4739 VGND.n317 VGND.t394 83.1719
R4740 VGND.n1210 VGND.n1206 78.6829
R4741 VGND.n1288 VGND.n1287 78.6829
R4742 VGND.n1313 VGND.n1312 78.6829
R4743 VGND.n1338 VGND.n1337 78.6829
R4744 VGND.n1363 VGND.n1362 78.6829
R4745 VGND.n1391 VGND.n1222 78.6829
R4746 VGND.n1249 VGND.n1248 78.6829
R4747 VGND.n1398 VGND.n1397 78.6829
R4748 VGND.n1018 VGND.n1017 78.6611
R4749 VGND.n1394 VGND.n545 77.9686
R4750 VGND.n1210 VGND.n1209 77.9299
R4751 VGND.n1287 VGND.n1285 77.9299
R4752 VGND.n1312 VGND.n1310 77.9299
R4753 VGND.n1337 VGND.n1335 77.9299
R4754 VGND.n1362 VGND.n1360 77.9299
R4755 VGND.n1391 VGND.n1390 77.9299
R4756 VGND.n1248 VGND.n1247 77.9299
R4757 VGND.n1397 VGND.n533 77.9299
R4758 VGND.n201 VGND.n200 75.905
R4759 VGND.n197 VGND.n196 75.905
R4760 VGND.n178 VGND.n177 75.905
R4761 VGND.n174 VGND.n173 75.905
R4762 VGND.n848 VGND.n847 75.905
R4763 VGND.n845 VGND.n844 75.905
R4764 VGND.n834 VGND.n833 75.905
R4765 VGND.n831 VGND.n830 75.905
R4766 VGND.n820 VGND.n819 75.905
R4767 VGND.n817 VGND.n816 75.905
R4768 VGND.n806 VGND.n805 75.905
R4769 VGND.n803 VGND.n802 75.905
R4770 VGND.n793 VGND.n792 75.905
R4771 VGND.n768 VGND.n767 75.905
R4772 VGND.n735 VGND.n734 75.905
R4773 VGND.n731 VGND.n730 75.905
R4774 VGND.n1018 VGND.n725 74.8287
R4775 VGND.n316 VGND.n315 73.3531
R4776 VGND.n1205 VGND.n1204 73.1255
R4777 VGND.n1204 VGND.n1168 73.1255
R4778 VGND.n1291 VGND.n1289 73.1255
R4779 VGND.n1291 VGND.n1168 73.1255
R4780 VGND.n1316 VGND.n1314 73.1255
R4781 VGND.n1316 VGND.n1168 73.1255
R4782 VGND.n1341 VGND.n1339 73.1255
R4783 VGND.n1341 VGND.n1168 73.1255
R4784 VGND.n1366 VGND.n1364 73.1255
R4785 VGND.n1366 VGND.n1168 73.1255
R4786 VGND.n1230 VGND.n1229 73.1255
R4787 VGND.n1230 VGND.n1168 73.1255
R4788 VGND.n1251 VGND.n1250 73.1255
R4789 VGND.n1251 VGND.n1168 73.1255
R4790 VGND.n1185 VGND.n554 73.1255
R4791 VGND.n1185 VGND.n1168 73.1255
R4792 VGND.n883 VGND.n850 73.1255
R4793 VGND.n850 VGND.n160 73.1255
R4794 VGND.n889 VGND.n887 73.1255
R4795 VGND.n887 VGND.n160 73.1255
R4796 VGND.n905 VGND.n836 73.1255
R4797 VGND.n836 VGND.n160 73.1255
R4798 VGND.n911 VGND.n909 73.1255
R4799 VGND.n909 VGND.n160 73.1255
R4800 VGND.n927 VGND.n822 73.1255
R4801 VGND.n822 VGND.n160 73.1255
R4802 VGND.n933 VGND.n931 73.1255
R4803 VGND.n931 VGND.n160 73.1255
R4804 VGND.n949 VGND.n808 73.1255
R4805 VGND.n808 VGND.n160 73.1255
R4806 VGND.n955 VGND.n953 73.1255
R4807 VGND.n953 VGND.n160 73.1255
R4808 VGND.n791 VGND.n790 73.1255
R4809 VGND.n790 VGND.n160 73.1255
R4810 VGND.n979 VGND.n770 73.1255
R4811 VGND.n770 VGND.n160 73.1255
R4812 VGND.n1008 VGND.n737 73.1255
R4813 VGND.n1002 VGND.n737 73.1255
R4814 VGND.n727 VGND.n726 73.1255
R4815 VGND.n997 VGND.n726 73.1255
R4816 VGND.n306 VGND.n190 73.1255
R4817 VGND.n313 VGND.n190 73.1255
R4818 VGND.n312 VGND.n311 73.1255
R4819 VGND.n313 VGND.n312 73.1255
R4820 VGND.n320 VGND.n180 73.1255
R4821 VGND.n187 VGND.n180 73.1255
R4822 VGND.n170 VGND.n169 73.1255
R4823 VGND.n182 VGND.n169 73.1255
R4824 VGND.n1712 VGND.t41 71.4713
R4825 VGND.n1752 VGND.n163 69.2272
R4826 VGND.n1756 VGND.n156 69.2272
R4827 VGND.n266 VGND.n265 69.2272
R4828 VGND.n232 VGND.n231 69.2272
R4829 VGND.n303 VGND.n191 68.7758
R4830 VGND.n299 VGND.n284 68.7561
R4831 VGND.n285 VGND.n284 68.7561
R4832 VGND.n292 VGND.n286 68.7561
R4833 VGND.n292 VGND.n291 68.7561
R4834 VGND.n280 VGND.n211 68.7561
R4835 VGND.n212 VGND.n211 68.7561
R4836 VGND.n273 VGND.n213 68.7561
R4837 VGND.n273 VGND.n272 68.7561
R4838 VGND.n244 VGND.n235 68.7561
R4839 VGND.n244 VGND.n243 68.7561
R4840 VGND.n993 VGND.n738 68.7561
R4841 VGND.n993 VGND.n992 68.7561
R4842 VGND.n987 VGND.n764 68.7561
R4843 VGND.n765 VGND.n764 68.7561
R4844 VGND.n966 VGND.n795 68.7561
R4845 VGND.n966 VGND.n965 68.7561
R4846 VGND.n961 VGND.n798 68.7561
R4847 VGND.n961 VGND.n960 68.7561
R4848 VGND.n944 VGND.n809 68.7561
R4849 VGND.n944 VGND.n943 68.7561
R4850 VGND.n939 VGND.n812 68.7561
R4851 VGND.n939 VGND.n938 68.7561
R4852 VGND.n922 VGND.n823 68.7561
R4853 VGND.n922 VGND.n921 68.7561
R4854 VGND.n917 VGND.n826 68.7561
R4855 VGND.n917 VGND.n916 68.7561
R4856 VGND.n900 VGND.n837 68.7561
R4857 VGND.n900 VGND.n899 68.7561
R4858 VGND.n895 VGND.n840 68.7561
R4859 VGND.n895 VGND.n894 68.7561
R4860 VGND.n878 VGND.n851 68.7561
R4861 VGND.n878 VGND.n877 68.7561
R4862 VGND.n873 VGND.n854 68.7561
R4863 VGND.n873 VGND.n872 68.7561
R4864 VGND.n1775 VGND.n1774 68.7561
R4865 VGND.n1789 VGND.n86 68.7561
R4866 VGND.n1806 VGND.n1805 68.7561
R4867 VGND.n511 VGND.n340 68.7561
R4868 VGND.n153 VGND.n144 68.7561
R4869 VGND.n149 VGND.n144 68.7561
R4870 VGND.t292 VGND.t474 68.6043
R4871 VGND.t18 VGND.t476 68.6043
R4872 VGND.t407 VGND.t482 68.6043
R4873 VGND.t399 VGND.t396 68.6043
R4874 VGND.n234 VGND.n233 67.5509
R4875 VGND.n218 VGND.n217 67.5509
R4876 VGND.n862 VGND.n861 67.5509
R4877 VGND.n860 VGND.n859 67.5509
R4878 VGND.n1734 VGND.n339 67.1161
R4879 VGND.n1046 VGND.n1044 67.1161
R4880 VGND.n1031 VGND.n1029 67.1161
R4881 VGND.n1059 VGND.n706 67.1161
R4882 VGND.n1062 VGND.n703 67.1161
R4883 VGND.n693 VGND.n692 67.1161
R4884 VGND.n691 VGND.n689 67.1161
R4885 VGND.n1085 VGND.n669 67.1161
R4886 VGND.n667 VGND.n665 67.1161
R4887 VGND.n1098 VGND.n645 67.1161
R4888 VGND.n643 VGND.n641 67.1161
R4889 VGND.n1111 VGND.n621 67.1161
R4890 VGND.n619 VGND.n617 67.1161
R4891 VGND.n1124 VGND.n597 67.1161
R4892 VGND.n595 VGND.n593 67.1161
R4893 VGND.n1137 VGND.n575 67.1161
R4894 VGND.n1800 VGND.n70 66.9639
R4895 VGND.n1799 VGND.n71 66.9639
R4896 VGND.n73 VGND.n72 66.9639
R4897 VGND.n1643 VGND.n1642 66.9639
R4898 VGND.n1641 VGND.n1640 66.9639
R4899 VGND.n1638 VGND.n1637 66.9639
R4900 VGND.n1661 VGND.n1636 66.9639
R4901 VGND.n1662 VGND.n1635 66.9639
R4902 VGND.n1665 VGND.n1632 66.9639
R4903 VGND.n1666 VGND.n1631 66.9639
R4904 VGND.n1668 VGND.n1630 66.9639
R4905 VGND.n1669 VGND.n1629 66.9639
R4906 VGND.n1617 VGND.n1616 66.9639
R4907 VGND.n1614 VGND.n1613 66.9639
R4908 VGND.n1679 VGND.n1612 66.9639
R4909 VGND.n1680 VGND.n1611 66.9639
R4910 VGND.n1683 VGND.n1608 66.9639
R4911 VGND.n1684 VGND.n1607 66.9639
R4912 VGND.n1686 VGND.n1606 66.9639
R4913 VGND.n1687 VGND.n1605 66.9639
R4914 VGND.n1593 VGND.n1592 66.9639
R4915 VGND.n1590 VGND.n1589 66.9639
R4916 VGND.n1697 VGND.n1588 66.9639
R4917 VGND.n1698 VGND.n1587 66.9639
R4918 VGND.n1701 VGND.n1584 66.9639
R4919 VGND.n1702 VGND.n1583 66.9639
R4920 VGND.n1704 VGND.n1582 66.9639
R4921 VGND.n1705 VGND.n1581 66.9639
R4922 VGND.n1529 VGND.n1528 66.9639
R4923 VGND.n1527 VGND.n1526 66.9639
R4924 VGND.n1540 VGND.n1525 66.9639
R4925 VGND.n1541 VGND.n1524 66.9639
R4926 VGND.n1522 VGND.n1403 66.9639
R4927 VGND.n1521 VGND.n1404 66.9639
R4928 VGND.n1519 VGND.n1405 66.9639
R4929 VGND.n1518 VGND.n1406 66.9639
R4930 VGND.n1515 VGND.n1413 66.9639
R4931 VGND.n1514 VGND.n1414 66.9639
R4932 VGND.n1416 VGND.n1415 66.9639
R4933 VGND.n1509 VGND.n1508 66.9639
R4934 VGND.n1506 VGND.n1425 66.9639
R4935 VGND.n1505 VGND.n1426 66.9639
R4936 VGND.n1428 VGND.n1427 66.9639
R4937 VGND.n1500 VGND.n1499 66.9639
R4938 VGND.n1497 VGND.n1437 66.9639
R4939 VGND.n1496 VGND.n1438 66.9639
R4940 VGND.n1440 VGND.n1439 66.9639
R4941 VGND.n1491 VGND.n1490 66.9639
R4942 VGND.n1488 VGND.n1449 66.9639
R4943 VGND.n1487 VGND.n1450 66.9639
R4944 VGND.n1452 VGND.n1451 66.9639
R4945 VGND.n1482 VGND.n1481 66.9639
R4946 VGND.n1479 VGND.n1461 66.9639
R4947 VGND.n1478 VGND.n1462 66.9639
R4948 VGND.n1464 VGND.n1463 66.9639
R4949 VGND.n1473 VGND.n1472 66.9639
R4950 VGND.n1157 VGND.n1156 66.9639
R4951 VGND.n1154 VGND.n1153 66.9639
R4952 VGND.n1555 VGND.n1152 66.9639
R4953 VGND.n1556 VGND.n1151 66.9639
R4954 VGND.n1559 VGND.n1144 66.9639
R4955 VGND.n1560 VGND.n1143 66.9639
R4956 VGND.n1562 VGND.n1142 66.9639
R4957 VGND.n1563 VGND.n1141 66.9639
R4958 VGND.n252 VGND.n227 65.0005
R4959 VGND.n259 VGND.n258 65.0005
R4960 VGND.n1760 VGND.n1759 65.0005
R4961 VGND.n165 VGND.n138 65.0005
R4962 VGND.n1758 VGND.n140 65.0005
R4963 VGND.n1748 VGND.n140 65.0005
R4964 VGND.n1750 VGND.n1749 65.0005
R4965 VGND.n1749 VGND.n1748 65.0005
R4966 VGND.n254 VGND.n253 65.0005
R4967 VGND.n255 VGND.n254 65.0005
R4968 VGND.n257 VGND.n256 65.0005
R4969 VGND.n256 VGND.n255 65.0005
R4970 VGND.n1019 VGND.t465 61.0779
R4971 VGND.n1041 VGND.t302 61.0779
R4972 VGND.n1713 VGND.t158 59.2465
R4973 VGND.n1026 VGND.t237 58.651
R4974 VGND.t194 VGND.n1026 58.651
R4975 VGND.t558 VGND.n1051 58.651
R4976 VGND.n1739 VGND.t341 58.651
R4977 VGND.t348 VGND.n1739 58.651
R4978 VGND.t97 VGND.n332 58.651
R4979 VGND.n1765 VGND.n1764 58.5005
R4980 VGND.n1764 VGND.n1763 58.5005
R4981 VGND.n1833 VGND.n3 58.5005
R4982 VGND.n239 VGND.n3 58.5005
R4983 VGND.n1754 VGND.n159 57.2454
R4984 VGND.n1713 VGND.t437 56.6133
R4985 VGND.n303 VGND.t26 55.8298
R4986 VGND.n1830 VGND.t294 55.0911
R4987 VGND.n1003 VGND.n135 53.6536
R4988 VGND.t502 VGND.t504 50.8275
R4989 VGND.t16 VGND.t542 50.8275
R4990 VGND.t403 VGND.t126 50.8275
R4991 VGND.t394 VGND.t405 50.8275
R4992 VGND.t200 VGND.n262 50.614
R4993 VGND.n1548 VGND.n1400 50.16
R4994 VGND.n1776 VGND.n125 49.4227
R4995 VGND.n1778 VGND.n119 49.4227
R4996 VGND.n1780 VGND.n113 49.4227
R4997 VGND.n1782 VGND.n107 49.4227
R4998 VGND.n1784 VGND.n101 49.4227
R4999 VGND.n1786 VGND.n95 49.4227
R5000 VGND.n1788 VGND.n89 49.4227
R5001 VGND.n1807 VGND.n63 49.4227
R5002 VGND.n1809 VGND.n57 49.4227
R5003 VGND.n1811 VGND.n51 49.4227
R5004 VGND.n1813 VGND.n45 49.4227
R5005 VGND.n1815 VGND.n39 49.4227
R5006 VGND.n1817 VGND.n33 49.4227
R5007 VGND.n1819 VGND.n27 49.4227
R5008 VGND.n1821 VGND.n21 49.4227
R5009 VGND.n471 VGND.n18 49.4227
R5010 VGND.n476 VGND.n467 49.4227
R5011 VGND.n478 VGND.n461 49.4227
R5012 VGND.n480 VGND.n455 49.4227
R5013 VGND.n482 VGND.n449 49.4227
R5014 VGND.n484 VGND.n443 49.4227
R5015 VGND.n486 VGND.n437 49.4227
R5016 VGND.n488 VGND.n431 49.4227
R5017 VGND.n490 VGND.n425 49.4227
R5018 VGND.n492 VGND.n419 49.4227
R5019 VGND.n494 VGND.n413 49.4227
R5020 VGND.n496 VGND.n407 49.4227
R5021 VGND.n498 VGND.n401 49.4227
R5022 VGND.n500 VGND.n395 49.4227
R5023 VGND.n502 VGND.n389 49.4227
R5024 VGND.n504 VGND.n383 49.4227
R5025 VGND.n506 VGND.n377 49.4227
R5026 VGND.n367 VGND.n365 49.4227
R5027 VGND.n369 VGND.n342 49.4227
R5028 VGND.n1726 VGND.n520 48.8605
R5029 VGND.t546 VGND.n1712 48.7138
R5030 VGND.n1743 VGND.n335 48.3561
R5031 VGND.n1737 VGND.n336 48.3561
R5032 VGND.n1043 VGND.n1032 48.3561
R5033 VGND.n1049 VGND.n710 48.3561
R5034 VGND.n1055 VGND.n709 48.3561
R5035 VGND.n714 VGND.n705 48.3561
R5036 VGND.n723 VGND.n704 48.3561
R5037 VGND.n702 VGND.n700 48.3561
R5038 VGND.n1075 VGND.n673 48.3561
R5039 VGND.n1081 VGND.n672 48.3561
R5040 VGND.n677 VGND.n668 48.3561
R5041 VGND.n1088 VGND.n649 48.3561
R5042 VGND.n1094 VGND.n648 48.3561
R5043 VGND.n653 VGND.n644 48.3561
R5044 VGND.n1101 VGND.n625 48.3561
R5045 VGND.n1107 VGND.n624 48.3561
R5046 VGND.n629 VGND.n620 48.3561
R5047 VGND.n1114 VGND.n601 48.3561
R5048 VGND.n1120 VGND.n600 48.3561
R5049 VGND.n605 VGND.n596 48.3561
R5050 VGND.n1127 VGND.n579 48.3561
R5051 VGND.n1133 VGND.n578 48.3561
R5052 VGND.n584 VGND.n574 48.3561
R5053 VGND.n1072 VGND.n694 48.3561
R5054 VGND.n1205 VGND.n1200 48.2672
R5055 VGND.n1295 VGND.n1289 48.2672
R5056 VGND.n1320 VGND.n1314 48.2672
R5057 VGND.n1345 VGND.n1339 48.2672
R5058 VGND.n1370 VGND.n1364 48.2672
R5059 VGND.n1229 VGND.n1228 48.2672
R5060 VGND.n1250 VGND.n1241 48.2672
R5061 VGND.n1716 VGND.n554 48.2672
R5062 VGND.n329 VGND.n168 46.7844
R5063 VGND.n1200 VGND.n1199 46.7472
R5064 VGND.n1296 VGND.n1295 46.7472
R5065 VGND.n1321 VGND.n1320 46.7472
R5066 VGND.n1346 VGND.n1345 46.7472
R5067 VGND.n1371 VGND.n1370 46.7472
R5068 VGND.n1228 VGND.n1227 46.7472
R5069 VGND.n1243 VGND.n1241 46.7472
R5070 VGND.n1717 VGND.n1716 46.7472
R5071 VGND.n1212 VGND.n1211 45.0005
R5072 VGND.n1394 VGND.n1212 45.0005
R5073 VGND.n1286 VGND.n1215 45.0005
R5074 VGND.n1394 VGND.n1215 45.0005
R5075 VGND.n1311 VGND.n1195 45.0005
R5076 VGND.n1394 VGND.n1195 45.0005
R5077 VGND.n1336 VGND.n1218 45.0005
R5078 VGND.n1394 VGND.n1218 45.0005
R5079 VGND.n1361 VGND.n1192 45.0005
R5080 VGND.n1394 VGND.n1192 45.0005
R5081 VGND.n1393 VGND.n1392 45.0005
R5082 VGND.n1394 VGND.n1393 45.0005
R5083 VGND.n1242 VGND.n1189 45.0005
R5084 VGND.n1394 VGND.n1189 45.0005
R5085 VGND.n1396 VGND.n1395 45.0005
R5086 VGND.n1395 VGND.n1394 45.0005
R5087 VGND.n1022 VGND.n1021 42.4907
R5088 VGND.n1027 VGND.n712 42.4907
R5089 VGND.n1035 VGND.n1033 42.4907
R5090 VGND.n1744 VGND.n333 42.4907
R5091 VGND.n586 VGND.n585 42.4907
R5092 VGND.n591 VGND.n581 42.4907
R5093 VGND.n610 VGND.n609 42.4907
R5094 VGND.n615 VGND.n603 42.4907
R5095 VGND.n634 VGND.n633 42.4907
R5096 VGND.n639 VGND.n627 42.4907
R5097 VGND.n658 VGND.n657 42.4907
R5098 VGND.n663 VGND.n651 42.4907
R5099 VGND.n682 VGND.n681 42.4907
R5100 VGND.n687 VGND.n675 42.4907
R5101 VGND.n697 VGND.n695 42.4907
R5102 VGND.n724 VGND.n717 42.4907
R5103 VGND.n2 VGND.t156 42.0841
R5104 VGND.n1767 VGND.t154 42.0841
R5105 VGND.n234 VGND.t495 41.3938
R5106 VGND.n218 VGND.t493 41.3938
R5107 VGND.n862 VGND.t492 41.3938
R5108 VGND.n860 VGND.t494 41.3938
R5109 VGND.n530 VGND.n528 39.0005
R5110 VGND.n565 VGND.n528 39.0005
R5111 VGND.n518 VGND.n517 39.0005
R5112 VGND.n524 VGND.n518 39.0005
R5113 VGND.n1290 VGND.n1277 39.0005
R5114 VGND.n1290 VGND.n524 39.0005
R5115 VGND.n1315 VGND.n1274 39.0005
R5116 VGND.n1315 VGND.n524 39.0005
R5117 VGND.n1340 VGND.n1271 39.0005
R5118 VGND.n1340 VGND.n524 39.0005
R5119 VGND.n1365 VGND.n1268 39.0005
R5120 VGND.n1365 VGND.n524 39.0005
R5121 VGND.n1234 VGND.n1226 39.0005
R5122 VGND.n1226 VGND.n524 39.0005
R5123 VGND.n1259 VGND.n1240 39.0005
R5124 VGND.n1240 VGND.n524 39.0005
R5125 VGND.n141 VGND.n139 39.0005
R5126 VGND.n781 VGND.n139 39.0005
R5127 VGND.n858 VGND.n857 39.0005
R5128 VGND.n857 VGND.n781 39.0005
R5129 VGND.n251 VGND.n226 39.0005
R5130 VGND.n261 VGND.n226 39.0005
R5131 VGND.n260 VGND.n216 39.0005
R5132 VGND.n261 VGND.n260 39.0005
R5133 VGND.n582 VGND.t167 38.0445
R5134 VGND.n607 VGND.t335 38.0445
R5135 VGND.n631 VGND.t417 38.0445
R5136 VGND.n655 VGND.t190 38.0445
R5137 VGND.n679 VGND.t174 38.0445
R5138 VGND.n1070 VGND.t208 38.0445
R5139 VGND.t146 VGND.n80 37.3437
R5140 VGND.n722 VGND.n721 36.563
R5141 VGND.n721 VGND.n720 36.563
R5142 VGND.n1068 VGND.n1067 36.563
R5143 VGND.n1069 VGND.n1068 36.563
R5144 VGND.n1080 VGND.n1079 36.563
R5145 VGND.n1079 VGND.n1078 36.563
R5146 VGND.n683 VGND.n671 36.563
R5147 VGND.n684 VGND.n683 36.563
R5148 VGND.n1093 VGND.n1092 36.563
R5149 VGND.n1092 VGND.n1091 36.563
R5150 VGND.n659 VGND.n647 36.563
R5151 VGND.n660 VGND.n659 36.563
R5152 VGND.n1106 VGND.n1105 36.563
R5153 VGND.n1105 VGND.n1104 36.563
R5154 VGND.n635 VGND.n623 36.563
R5155 VGND.n636 VGND.n635 36.563
R5156 VGND.n1119 VGND.n1118 36.563
R5157 VGND.n1118 VGND.n1117 36.563
R5158 VGND.n611 VGND.n599 36.563
R5159 VGND.n612 VGND.n611 36.563
R5160 VGND.n1132 VGND.n1131 36.563
R5161 VGND.n1131 VGND.n1130 36.563
R5162 VGND.n587 VGND.n577 36.563
R5163 VGND.n588 VGND.n587 36.563
R5164 VGND.n1742 VGND.n1741 36.563
R5165 VGND.n1741 VGND.n1740 36.563
R5166 VGND.n1039 VGND.n1038 36.563
R5167 VGND.n1040 VGND.n1039 36.563
R5168 VGND.n1054 VGND.n1053 36.563
R5169 VGND.n1053 VGND.n1052 36.563
R5170 VGND.n1023 VGND.n708 36.563
R5171 VGND.n1024 VGND.n1023 36.563
R5172 VGND.n590 VGND.t201 36.5328
R5173 VGND.t35 VGND.n590 36.5328
R5174 VGND.t451 VGND.n1129 36.5328
R5175 VGND.n614 VGND.t459 36.5328
R5176 VGND.t470 VGND.n614 36.5328
R5177 VGND.t346 VGND.n1116 36.5328
R5178 VGND.n638 VGND.t256 36.5328
R5179 VGND.t7 VGND.n638 36.5328
R5180 VGND.t170 VGND.n1103 36.5328
R5181 VGND.n662 VGND.t483 36.5328
R5182 VGND.t532 VGND.n662 36.5328
R5183 VGND.t114 VGND.n1090 36.5328
R5184 VGND.n686 VGND.t339 36.5328
R5185 VGND.t13 VGND.n686 36.5328
R5186 VGND.t286 VGND.n1077 36.5328
R5187 VGND.n719 VGND.t95 36.5328
R5188 VGND.t128 VGND.n719 36.5328
R5189 VGND.t498 VGND.n715 36.5328
R5190 VGND.n1208 VGND.n1207 36.4805
R5191 VGND.n1299 VGND.n1298 36.4805
R5192 VGND.n1324 VGND.n1323 36.4805
R5193 VGND.n1349 VGND.n1348 36.4805
R5194 VGND.n1374 VGND.n1373 36.4805
R5195 VGND.n1389 VGND.n1388 36.4805
R5196 VGND.n1246 VGND.n1245 36.4805
R5197 VGND.n1722 VGND.n1721 36.4805
R5198 VGND.t504 VGND.n168 36.388
R5199 VGND.n1719 VGND.n537 35.6059
R5200 VGND.t465 VGND.t92 35.5953
R5201 VGND.t237 VGND.t557 35.5953
R5202 VGND.t467 VGND.t194 35.5953
R5203 VGND.t42 VGND.t558 35.5953
R5204 VGND.t302 VGND.t411 35.5953
R5205 VGND.t555 VGND.t341 35.5953
R5206 VGND.t253 VGND.t348 35.5953
R5207 VGND.t2 VGND.t97 35.5953
R5208 VGND.n1199 VGND.n1198 35.2005
R5209 VGND.n1297 VGND.n1296 35.2005
R5210 VGND.n1322 VGND.n1321 35.2005
R5211 VGND.n1347 VGND.n1346 35.2005
R5212 VGND.n1372 VGND.n1371 35.2005
R5213 VGND.n1227 VGND.n1221 35.2005
R5214 VGND.n1244 VGND.n1243 35.2005
R5215 VGND.n1717 VGND.n534 35.2005
R5216 VGND.n1038 VGND.n1032 35.1378
R5217 VGND.n714 VGND.n708 35.1378
R5218 VGND.n677 VGND.n671 35.1378
R5219 VGND.n653 VGND.n647 35.1378
R5220 VGND.n629 VGND.n623 35.1378
R5221 VGND.n605 VGND.n599 35.1378
R5222 VGND.n584 VGND.n577 35.1378
R5223 VGND.n1067 VGND.n694 35.1378
R5224 VGND.n1038 VGND.n1037 34.7613
R5225 VGND.n1742 VGND.n336 34.7613
R5226 VGND.n1743 VGND.n1742 34.7613
R5227 VGND.n1056 VGND.n708 34.7613
R5228 VGND.n1055 VGND.n1054 34.7613
R5229 VGND.n1054 VGND.n710 34.7613
R5230 VGND.n1082 VGND.n671 34.7613
R5231 VGND.n1081 VGND.n1080 34.7613
R5232 VGND.n1080 VGND.n673 34.7613
R5233 VGND.n1095 VGND.n647 34.7613
R5234 VGND.n1094 VGND.n1093 34.7613
R5235 VGND.n1093 VGND.n649 34.7613
R5236 VGND.n1108 VGND.n623 34.7613
R5237 VGND.n1107 VGND.n1106 34.7613
R5238 VGND.n1106 VGND.n625 34.7613
R5239 VGND.n1121 VGND.n599 34.7613
R5240 VGND.n1120 VGND.n1119 34.7613
R5241 VGND.n1119 VGND.n601 34.7613
R5242 VGND.n1134 VGND.n577 34.7613
R5243 VGND.n1133 VGND.n1132 34.7613
R5244 VGND.n1132 VGND.n579 34.7613
R5245 VGND.n1067 VGND.n1066 34.7613
R5246 VGND.n722 VGND.n700 34.7613
R5247 VGND.n723 VGND.n722 34.7613
R5248 VGND.n997 VGND.t292 34.3024
R5249 VGND.t476 VGND.n997 34.3024
R5250 VGND.n1002 VGND.t407 34.3024
R5251 VGND.t396 VGND.n1002 34.3024
R5252 VGND.n1207 VGND.n1198 32.9605
R5253 VGND.n1298 VGND.n1297 32.9605
R5254 VGND.n1323 VGND.n1322 32.9605
R5255 VGND.n1348 VGND.n1347 32.9605
R5256 VGND.n1373 VGND.n1372 32.9605
R5257 VGND.n1388 VGND.n1221 32.9605
R5258 VGND.n1245 VGND.n1244 32.9605
R5259 VGND.n1721 VGND.n534 32.9605
R5260 VGND.n1282 VGND.t162 31.7728
R5261 VGND.n1307 VGND.t457 31.7728
R5262 VGND.n1332 VGND.t145 31.7728
R5263 VGND.n1357 VGND.t435 31.7728
R5264 VGND.n1382 VGND.t228 31.7728
R5265 VGND.n1264 VGND.t458 31.7728
R5266 VGND.n1257 VGND.t116 31.7728
R5267 VGND.n572 VGND.t159 31.7728
R5268 VGND.n1748 VGND.t124 31.6536
R5269 VGND.n1034 VGND.n166 31.1459
R5270 VGND.n330 VGND.n329 30.6122
R5271 VGND.n1407 VGND.n1402 28.8579
R5272 VGND.n1512 VGND.n1417 28.8579
R5273 VGND.n1503 VGND.n1429 28.8579
R5274 VGND.n1494 VGND.n1441 28.8579
R5275 VGND.n1485 VGND.n1453 28.8579
R5276 VGND.n1476 VGND.n1465 28.8579
R5277 VGND.n1553 VGND.n1155 28.8579
R5278 VGND.n1145 VGND.n567 28.8579
R5279 VGND.n1659 VGND.n1639 28.8579
R5280 VGND.n1647 VGND.n1628 28.8579
R5281 VGND.n1677 VGND.n1615 28.8579
R5282 VGND.n1620 VGND.n1604 28.8579
R5283 VGND.n1695 VGND.n1591 28.8579
R5284 VGND.n1596 VGND.n1580 28.8579
R5285 VGND.n1538 VGND.n1537 28.857
R5286 VGND.n1797 VGND.n1796 28.857
R5287 VGND.n1537 VGND.n1536 28.6936
R5288 VGND.n1796 VGND.n1795 28.6936
R5289 VGND.n1597 VGND.n1596 28.6927
R5290 VGND.n1602 VGND.n1591 28.6927
R5291 VGND.n1621 VGND.n1620 28.6927
R5292 VGND.n1626 VGND.n1615 28.6927
R5293 VGND.n1648 VGND.n1647 28.6927
R5294 VGND.n1653 VGND.n1639 28.6927
R5295 VGND.n1146 VGND.n1145 28.6927
R5296 VGND.n1162 VGND.n1155 28.6927
R5297 VGND.n1469 VGND.n1465 28.6927
R5298 VGND.n1457 VGND.n1453 28.6927
R5299 VGND.n1445 VGND.n1441 28.6927
R5300 VGND.n1433 VGND.n1429 28.6927
R5301 VGND.n1421 VGND.n1417 28.6927
R5302 VGND.n1408 VGND.n1407 28.6927
R5303 VGND.n1746 VGND.n1745 28.3145
R5304 VGND.t26 VGND.n301 26.7015
R5305 VGND.t491 VGND.n160 26.0413
R5306 VGND.n516 VGND.n515 25.9728
R5307 VGND.n1281 VGND.n1280 25.9728
R5308 VGND.n1305 VGND.n1279 25.9728
R5309 VGND.n1306 VGND.n1278 25.9728
R5310 VGND.n1330 VGND.n1276 25.9728
R5311 VGND.n1331 VGND.n1275 25.9728
R5312 VGND.n1355 VGND.n1273 25.9728
R5313 VGND.n1356 VGND.n1272 25.9728
R5314 VGND.n1380 VGND.n1270 25.9728
R5315 VGND.n1381 VGND.n1269 25.9728
R5316 VGND.n1266 VGND.n1224 25.9728
R5317 VGND.n1265 VGND.n1225 25.9728
R5318 VGND.n1239 VGND.n1238 25.9728
R5319 VGND.n1256 VGND.n1255 25.9728
R5320 VGND.n570 VGND.n569 25.9728
R5321 VGND.n571 VGND.n568 25.9728
R5322 VGND.n1733 VGND.n335 25.8532
R5323 VGND.n1737 VGND.n1736 25.8532
R5324 VGND.n1047 VGND.n1043 25.8532
R5325 VGND.n1049 VGND.n1048 25.8532
R5326 VGND.n709 VGND.n707 25.8532
R5327 VGND.n1060 VGND.n705 25.8532
R5328 VGND.n1061 VGND.n704 25.8532
R5329 VGND.n1064 VGND.n702 25.8532
R5330 VGND.n1075 VGND.n1074 25.8532
R5331 VGND.n672 VGND.n670 25.8532
R5332 VGND.n1086 VGND.n668 25.8532
R5333 VGND.n1088 VGND.n1087 25.8532
R5334 VGND.n648 VGND.n646 25.8532
R5335 VGND.n1099 VGND.n644 25.8532
R5336 VGND.n1101 VGND.n1100 25.8532
R5337 VGND.n624 VGND.n622 25.8532
R5338 VGND.n1112 VGND.n620 25.8532
R5339 VGND.n1114 VGND.n1113 25.8532
R5340 VGND.n600 VGND.n598 25.8532
R5341 VGND.n1125 VGND.n596 25.8532
R5342 VGND.n1127 VGND.n1126 25.8532
R5343 VGND.n578 VGND.n576 25.8532
R5344 VGND.n1138 VGND.n574 25.8532
R5345 VGND.n1073 VGND.n1072 25.8532
R5346 VGND.n182 VGND.t502 25.414
R5347 VGND.t542 VGND.n182 25.414
R5348 VGND.n187 VGND.t403 25.414
R5349 VGND.t405 VGND.n187 25.414
R5350 VGND.n157 VGND.n156 24.3755
R5351 VGND.n159 VGND.n157 24.3755
R5352 VGND.n163 VGND.n161 24.3755
R5353 VGND.n161 VGND.n159 24.3755
R5354 VGND.n232 VGND.n230 24.3755
R5355 VGND.n230 VGND.n189 24.3755
R5356 VGND.n266 VGND.n220 24.3755
R5357 VGND.n220 VGND.n189 24.3755
R5358 VGND.n1201 VGND.n1200 23.1494
R5359 VGND.n1295 VGND.n1294 23.1494
R5360 VGND.n1320 VGND.n1319 23.1494
R5361 VGND.n1345 VGND.n1344 23.1494
R5362 VGND.n1370 VGND.n1369 23.1494
R5363 VGND.n1233 VGND.n1228 23.1494
R5364 VGND.n1254 VGND.n1241 23.1494
R5365 VGND.n1716 VGND.n1715 23.1494
R5366 VGND.n1719 VGND.n545 23.131
R5367 VGND.n1302 VGND.n1301 22.5005
R5368 VGND.n1301 VGND.n537 22.5005
R5369 VGND.n1327 VGND.n1326 22.5005
R5370 VGND.n1326 VGND.n537 22.5005
R5371 VGND.n1352 VGND.n1351 22.5005
R5372 VGND.n1351 VGND.n537 22.5005
R5373 VGND.n1377 VGND.n1376 22.5005
R5374 VGND.n1376 VGND.n537 22.5005
R5375 VGND.n1387 VGND.n1386 22.5005
R5376 VGND.n1386 VGND.n537 22.5005
R5377 VGND.n1237 VGND.n1236 22.5005
R5378 VGND.n1236 VGND.n537 22.5005
R5379 VGND.n1723 VGND.n529 22.5005
R5380 VGND.n537 VGND.n529 22.5005
R5381 VGND.n519 VGND.n514 22.5005
R5382 VGND.n1711 VGND.n519 22.5005
R5383 VGND.t167 VGND.t37 22.1718
R5384 VGND.t201 VGND.t157 22.1718
R5385 VGND.t169 VGND.t35 22.1718
R5386 VGND.t119 VGND.t451 22.1718
R5387 VGND.t335 VGND.t496 22.1718
R5388 VGND.t459 VGND.t345 22.1718
R5389 VGND.t334 VGND.t470 22.1718
R5390 VGND.t225 VGND.t346 22.1718
R5391 VGND.t417 VGND.t245 22.1718
R5392 VGND.t256 VGND.t107 22.1718
R5393 VGND.t99 VGND.t7 22.1718
R5394 VGND.t472 VGND.t170 22.1718
R5395 VGND.t190 VGND.t242 22.1718
R5396 VGND.t483 VGND.t221 22.1718
R5397 VGND.t365 VGND.t532 22.1718
R5398 VGND.t32 VGND.t114 22.1718
R5399 VGND.t174 VGND.t87 22.1718
R5400 VGND.t339 VGND.t140 22.1718
R5401 VGND.t311 VGND.t13 22.1718
R5402 VGND.t552 VGND.t286 22.1718
R5403 VGND.t208 VGND.t117 22.1718
R5404 VGND.t95 VGND.t210 22.1718
R5405 VGND.t283 VGND.t128 22.1718
R5406 VGND.t550 VGND.t498 22.1718
R5407 VGND.t41 VGND.n524 20.0123
R5408 VGND.n1712 VGND.n1711 19.4911
R5409 VGND.n1789 VGND.n1788 19.3338
R5410 VGND.n1788 VGND.n1787 19.3338
R5411 VGND.n1787 VGND.n1786 19.3338
R5412 VGND.n1786 VGND.n1785 19.3338
R5413 VGND.n1785 VGND.n1784 19.3338
R5414 VGND.n1784 VGND.n1783 19.3338
R5415 VGND.n1783 VGND.n1782 19.3338
R5416 VGND.n1782 VGND.n1781 19.3338
R5417 VGND.n1781 VGND.n1780 19.3338
R5418 VGND.n1780 VGND.n1779 19.3338
R5419 VGND.n1779 VGND.n1778 19.3338
R5420 VGND.n1778 VGND.n1777 19.3338
R5421 VGND.n1777 VGND.n1776 19.3338
R5422 VGND.n1776 VGND.n1775 19.3338
R5423 VGND.n511 VGND.n342 19.3338
R5424 VGND.n371 VGND.n342 19.3338
R5425 VGND.n371 VGND.n365 19.3338
R5426 VGND.n507 VGND.n365 19.3338
R5427 VGND.n507 VGND.n506 19.3338
R5428 VGND.n506 VGND.n505 19.3338
R5429 VGND.n505 VGND.n504 19.3338
R5430 VGND.n504 VGND.n503 19.3338
R5431 VGND.n503 VGND.n502 19.3338
R5432 VGND.n502 VGND.n501 19.3338
R5433 VGND.n501 VGND.n500 19.3338
R5434 VGND.n500 VGND.n499 19.3338
R5435 VGND.n499 VGND.n498 19.3338
R5436 VGND.n498 VGND.n497 19.3338
R5437 VGND.n497 VGND.n496 19.3338
R5438 VGND.n496 VGND.n495 19.3338
R5439 VGND.n495 VGND.n494 19.3338
R5440 VGND.n494 VGND.n493 19.3338
R5441 VGND.n493 VGND.n492 19.3338
R5442 VGND.n492 VGND.n491 19.3338
R5443 VGND.n491 VGND.n490 19.3338
R5444 VGND.n490 VGND.n489 19.3338
R5445 VGND.n489 VGND.n488 19.3338
R5446 VGND.n488 VGND.n487 19.3338
R5447 VGND.n487 VGND.n486 19.3338
R5448 VGND.n486 VGND.n485 19.3338
R5449 VGND.n485 VGND.n484 19.3338
R5450 VGND.n484 VGND.n483 19.3338
R5451 VGND.n483 VGND.n482 19.3338
R5452 VGND.n482 VGND.n481 19.3338
R5453 VGND.n481 VGND.n480 19.3338
R5454 VGND.n480 VGND.n479 19.3338
R5455 VGND.n479 VGND.n478 19.3338
R5456 VGND.n478 VGND.n477 19.3338
R5457 VGND.n477 VGND.n476 19.3338
R5458 VGND.n476 VGND.n475 19.3338
R5459 VGND.n475 VGND.n18 19.3338
R5460 VGND.n1822 VGND.n18 19.3338
R5461 VGND.n1822 VGND.n1821 19.3338
R5462 VGND.n1821 VGND.n1820 19.3338
R5463 VGND.n1820 VGND.n1819 19.3338
R5464 VGND.n1819 VGND.n1818 19.3338
R5465 VGND.n1818 VGND.n1817 19.3338
R5466 VGND.n1817 VGND.n1816 19.3338
R5467 VGND.n1816 VGND.n1815 19.3338
R5468 VGND.n1815 VGND.n1814 19.3338
R5469 VGND.n1814 VGND.n1813 19.3338
R5470 VGND.n1813 VGND.n1812 19.3338
R5471 VGND.n1812 VGND.n1811 19.3338
R5472 VGND.n1811 VGND.n1810 19.3338
R5473 VGND.n1810 VGND.n1809 19.3338
R5474 VGND.n1809 VGND.n1808 19.3338
R5475 VGND.n1808 VGND.n1807 19.3338
R5476 VGND.n1807 VGND.n1806 19.3338
R5477 VGND.n976 VGND.n771 19.0821
R5478 VGND.t557 VGND.n1024 19.0113
R5479 VGND.n1040 VGND.t555 19.0113
R5480 VGND.n301 VGND.t74 18.6103
R5481 VGND.n1208 VGND.n514 18.2672
R5482 VGND.n1302 VGND.n1299 18.2672
R5483 VGND.n1327 VGND.n1324 18.2672
R5484 VGND.n1352 VGND.n1349 18.2672
R5485 VGND.n1377 VGND.n1374 18.2672
R5486 VGND.n1389 VGND.n1387 18.2672
R5487 VGND.n1246 VGND.n1237 18.2672
R5488 VGND.n1723 VGND.n1722 18.2672
R5489 VGND.n354 VGND.t105 18.0461
R5490 VGND.n1052 VGND.t467 17.7979
R5491 VGND.n1052 VGND.t42 17.7979
R5492 VGND.n1740 VGND.t253 17.7979
R5493 VGND.n1740 VGND.t2 17.7979
R5494 VGND.n233 VGND.t416 17.4005
R5495 VGND.n233 VGND.t31 17.4005
R5496 VGND.n217 VGND.t83 17.4005
R5497 VGND.n217 VGND.t537 17.4005
R5498 VGND.n200 VGND.t398 17.4005
R5499 VGND.n200 VGND.t401 17.4005
R5500 VGND.n196 VGND.t27 17.4005
R5501 VGND.n196 VGND.t100 17.4005
R5502 VGND.n177 VGND.t404 17.4005
R5503 VGND.n177 VGND.t406 17.4005
R5504 VGND.n173 VGND.t503 17.4005
R5505 VGND.n173 VGND.t543 17.4005
R5506 VGND.n861 VGND.t166 17.4005
R5507 VGND.n861 VGND.t1 17.4005
R5508 VGND.n859 VGND.t207 17.4005
R5509 VGND.n859 VGND.t25 17.4005
R5510 VGND.n847 VGND.t299 17.4005
R5511 VGND.n847 VGND.t308 17.4005
R5512 VGND.n844 VGND.t529 17.4005
R5513 VGND.n844 VGND.t285 17.4005
R5514 VGND.n833 VGND.t151 17.4005
R5515 VGND.n833 VGND.t152 17.4005
R5516 VGND.n830 VGND.t359 17.4005
R5517 VGND.n830 VGND.t357 17.4005
R5518 VGND.n819 VGND.t186 17.4005
R5519 VGND.n819 VGND.t185 17.4005
R5520 VGND.n816 VGND.t143 17.4005
R5521 VGND.n816 VGND.t260 17.4005
R5522 VGND.n805 VGND.t361 17.4005
R5523 VGND.n805 VGND.t360 17.4005
R5524 VGND.n802 VGND.t291 17.4005
R5525 VGND.n802 VGND.t290 17.4005
R5526 VGND.n792 VGND.t91 17.4005
R5527 VGND.n792 VGND.t34 17.4005
R5528 VGND.n767 VGND.t203 17.4005
R5529 VGND.n767 VGND.t193 17.4005
R5530 VGND.n734 VGND.t408 17.4005
R5531 VGND.n734 VGND.t397 17.4005
R5532 VGND.n730 VGND.t293 17.4005
R5533 VGND.n730 VGND.t477 17.4005
R5534 VGND.n70 VGND.t371 17.4005
R5535 VGND.n70 VGND.t373 17.4005
R5536 VGND.n71 VGND.t367 17.4005
R5537 VGND.n71 VGND.t369 17.4005
R5538 VGND.n72 VGND.t381 17.4005
R5539 VGND.n72 VGND.t375 17.4005
R5540 VGND.n1642 VGND.t384 17.4005
R5541 VGND.n1642 VGND.t378 17.4005
R5542 VGND.n1640 VGND.t275 17.4005
R5543 VGND.n1640 VGND.t331 17.4005
R5544 VGND.n1637 VGND.t329 17.4005
R5545 VGND.n1637 VGND.t277 17.4005
R5546 VGND.n1636 VGND.t47 17.4005
R5547 VGND.n1636 VGND.t69 17.4005
R5548 VGND.n1635 VGND.t122 17.4005
R5549 VGND.n1635 VGND.t319 17.4005
R5550 VGND.n1632 VGND.t322 17.4005
R5551 VGND.n1632 VGND.t455 17.4005
R5552 VGND.n1631 VGND.t57 17.4005
R5553 VGND.n1631 VGND.t480 17.4005
R5554 VGND.n1630 VGND.t255 17.4005
R5555 VGND.n1630 VGND.t545 17.4005
R5556 VGND.n1629 VGND.t252 17.4005
R5557 VGND.n1629 VGND.t301 17.4005
R5558 VGND.n1616 VGND.t430 17.4005
R5559 VGND.n1616 VGND.t333 17.4005
R5560 VGND.n1613 VGND.t279 17.4005
R5561 VGND.n1613 VGND.t432 17.4005
R5562 VGND.n1612 VGND.t197 17.4005
R5563 VGND.n1612 VGND.t102 17.4005
R5564 VGND.n1611 VGND.t179 17.4005
R5565 VGND.n1611 VGND.t104 17.4005
R5566 VGND.n1608 VGND.t113 17.4005
R5567 VGND.n1608 VGND.t507 17.4005
R5568 VGND.n1607 VGND.t142 17.4005
R5569 VGND.n1607 VGND.t139 17.4005
R5570 VGND.n1606 VGND.t305 17.4005
R5571 VGND.n1606 VGND.t428 17.4005
R5572 VGND.n1605 VGND.t307 17.4005
R5573 VGND.n1605 VGND.t420 17.4005
R5574 VGND.n1592 VGND.t501 17.4005
R5575 VGND.n1592 VGND.t216 17.4005
R5576 VGND.n1589 VGND.t71 17.4005
R5577 VGND.n1589 VGND.t109 17.4005
R5578 VGND.n1588 VGND.t232 17.4005
R5579 VGND.n1588 VGND.t250 17.4005
R5580 VGND.n1587 VGND.t248 17.4005
R5581 VGND.n1587 VGND.t67 17.4005
R5582 VGND.n1584 VGND.t206 17.4005
R5583 VGND.n1584 VGND.t536 17.4005
R5584 VGND.n1583 VGND.t173 17.4005
R5585 VGND.n1583 VGND.t464 17.4005
R5586 VGND.n1582 VGND.t22 17.4005
R5587 VGND.n1582 VGND.t273 17.4005
R5588 VGND.n1581 VGND.t271 17.4005
R5589 VGND.n1581 VGND.t24 17.4005
R5590 VGND.n339 VGND.t3 17.4005
R5591 VGND.n339 VGND.t98 17.4005
R5592 VGND.n1044 VGND.t303 17.4005
R5593 VGND.n1044 VGND.t412 17.4005
R5594 VGND.n1029 VGND.t43 17.4005
R5595 VGND.n1029 VGND.t559 17.4005
R5596 VGND.n706 VGND.t466 17.4005
R5597 VGND.n706 VGND.t93 17.4005
R5598 VGND.n703 VGND.t551 17.4005
R5599 VGND.n703 VGND.t499 17.4005
R5600 VGND.n692 VGND.t209 17.4005
R5601 VGND.n692 VGND.t118 17.4005
R5602 VGND.n689 VGND.t553 17.4005
R5603 VGND.n689 VGND.t287 17.4005
R5604 VGND.n669 VGND.t175 17.4005
R5605 VGND.n669 VGND.t88 17.4005
R5606 VGND.n665 VGND.t33 17.4005
R5607 VGND.n665 VGND.t115 17.4005
R5608 VGND.n645 VGND.t191 17.4005
R5609 VGND.n645 VGND.t243 17.4005
R5610 VGND.n641 VGND.t473 17.4005
R5611 VGND.n641 VGND.t171 17.4005
R5612 VGND.n621 VGND.t418 17.4005
R5613 VGND.n621 VGND.t246 17.4005
R5614 VGND.n617 VGND.t226 17.4005
R5615 VGND.n617 VGND.t347 17.4005
R5616 VGND.n597 VGND.t336 17.4005
R5617 VGND.n597 VGND.t497 17.4005
R5618 VGND.n593 VGND.t120 17.4005
R5619 VGND.n593 VGND.t452 17.4005
R5620 VGND.n575 VGND.t168 17.4005
R5621 VGND.n575 VGND.t38 17.4005
R5622 VGND.n1528 VGND.t364 17.4005
R5623 VGND.n1528 VGND.t189 17.4005
R5624 VGND.n1526 VGND.t63 17.4005
R5625 VGND.n1526 VGND.t82 17.4005
R5626 VGND.n1525 VGND.t6 17.4005
R5627 VGND.n1525 VGND.t12 17.4005
R5628 VGND.n1524 VGND.t10 17.4005
R5629 VGND.n1524 VGND.t20 17.4005
R5630 VGND.n1403 VGND.t55 17.4005
R5631 VGND.n1403 VGND.t59 17.4005
R5632 VGND.n1404 VGND.t489 17.4005
R5633 VGND.n1404 VGND.t469 17.4005
R5634 VGND.n1405 VGND.t240 17.4005
R5635 VGND.n1405 VGND.t218 17.4005
R5636 VGND.n1406 VGND.t214 17.4005
R5637 VGND.n1406 VGND.t49 17.4005
R5638 VGND.n1413 VGND.t40 17.4005
R5639 VGND.n1413 VGND.t517 17.4005
R5640 VGND.n1414 VGND.t515 17.4005
R5641 VGND.n1414 VGND.t487 17.4005
R5642 VGND.n1415 VGND.t80 17.4005
R5643 VGND.n1415 VGND.t78 17.4005
R5644 VGND.n1508 VGND.t65 17.4005
R5645 VGND.n1508 VGND.t111 17.4005
R5646 VGND.n1425 VGND.t351 17.4005
R5647 VGND.n1425 VGND.t509 17.4005
R5648 VGND.n1426 VGND.t220 17.4005
R5649 VGND.n1426 VGND.t511 17.4005
R5650 VGND.n1427 VGND.t267 17.4005
R5651 VGND.n1427 VGND.t269 17.4005
R5652 VGND.n1499 VGND.t263 17.4005
R5653 VGND.n1499 VGND.t265 17.4005
R5654 VGND.n1437 VGND.t388 17.4005
R5655 VGND.n1437 VGND.t390 17.4005
R5656 VGND.n1438 VGND.t392 17.4005
R5657 VGND.n1438 VGND.t386 17.4005
R5658 VGND.n1439 VGND.t177 17.4005
R5659 VGND.n1439 VGND.t259 17.4005
R5660 VGND.n1490 VGND.t51 17.4005
R5661 VGND.n1490 VGND.t353 17.4005
R5662 VGND.n1449 VGND.t424 17.4005
R5663 VGND.n1449 VGND.t422 17.4005
R5664 VGND.n1450 VGND.t462 17.4005
R5665 VGND.n1450 VGND.t85 17.4005
R5666 VGND.n1451 VGND.t73 17.4005
R5667 VGND.n1451 VGND.t317 17.4005
R5668 VGND.n1481 VGND.t90 17.4005
R5669 VGND.n1481 VGND.t315 17.4005
R5670 VGND.n1461 VGND.t448 17.4005
R5671 VGND.n1461 VGND.t234 17.4005
R5672 VGND.n1462 VGND.t434 17.4005
R5673 VGND.n1462 VGND.t450 17.4005
R5674 VGND.n1463 VGND.t53 17.4005
R5675 VGND.n1463 VGND.t184 17.4005
R5676 VGND.n1472 VGND.t182 17.4005
R5677 VGND.n1472 VGND.t324 17.4005
R5678 VGND.n1156 VGND.t313 17.4005
R5679 VGND.n1156 VGND.t310 17.4005
R5680 VGND.n1153 VGND.t541 17.4005
R5681 VGND.n1153 VGND.t539 17.4005
R5682 VGND.n1152 VGND.t61 17.4005
R5683 VGND.n1152 VGND.t519 17.4005
R5684 VGND.n1151 VGND.t521 17.4005
R5685 VGND.n1151 VGND.t523 17.4005
R5686 VGND.n1144 VGND.t165 17.4005
R5687 VGND.n1144 VGND.t282 17.4005
R5688 VGND.n1143 VGND.t531 17.4005
R5689 VGND.n1143 VGND.t45 17.4005
R5690 VGND.n1142 VGND.t212 17.4005
R5691 VGND.n1142 VGND.t415 17.4005
R5692 VGND.n1141 VGND.t344 17.4005
R5693 VGND.n1141 VGND.t289 17.4005
R5694 VGND.n1762 VGND.t153 17.1575
R5695 VGND.n241 VGND.t294 16.6727
R5696 VGND.n1024 VGND.t92 16.5844
R5697 VGND.t411 VGND.n1040 16.5844
R5698 VGND.n1830 VGND.t155 15.9478
R5699 VGND.n1728 VGND.n1727 15.3952
R5700 VGND.n1727 VGND.n1726 15.3952
R5701 VGND.n1303 VGND.n525 15.3952
R5702 VGND.n1726 VGND.n525 15.3952
R5703 VGND.n1328 VGND.n523 15.3952
R5704 VGND.n1726 VGND.n523 15.3952
R5705 VGND.n1353 VGND.n526 15.3952
R5706 VGND.n1726 VGND.n526 15.3952
R5707 VGND.n1378 VGND.n522 15.3952
R5708 VGND.n1726 VGND.n522 15.3952
R5709 VGND.n1223 VGND.n527 15.3952
R5710 VGND.n1726 VGND.n527 15.3952
R5711 VGND.n1260 VGND.n521 15.3952
R5712 VGND.n1726 VGND.n521 15.3952
R5713 VGND.n1725 VGND.n1724 15.3952
R5714 VGND.n1726 VGND.n1725 15.3952
R5715 VGND.n976 VGND.n781 15.2658
R5716 VGND.t28 VGND.n11 14.0522
R5717 VGND.n1754 VGND.n160 11.8985
R5718 VGND.t157 VGND.n588 11.842
R5719 VGND.t345 VGND.n612 11.842
R5720 VGND.t107 VGND.n636 11.842
R5721 VGND.t221 VGND.n660 11.842
R5722 VGND.t140 VGND.n684 11.842
R5723 VGND.n1069 VGND.t210 11.842
R5724 VGND.n1130 VGND.t169 11.0862
R5725 VGND.n1130 VGND.t119 11.0862
R5726 VGND.n1117 VGND.t334 11.0862
R5727 VGND.n1117 VGND.t225 11.0862
R5728 VGND.n1104 VGND.t99 11.0862
R5729 VGND.n1104 VGND.t472 11.0862
R5730 VGND.n1091 VGND.t365 11.0862
R5731 VGND.n1091 VGND.t32 11.0862
R5732 VGND.n1078 VGND.t311 11.0862
R5733 VGND.n1078 VGND.t552 11.0862
R5734 VGND.n720 VGND.t283 11.0862
R5735 VGND.n720 VGND.t550 11.0862
R5736 VGND.n1394 VGND.t76 10.6561
R5737 VGND.n588 VGND.t37 10.3303
R5738 VGND.n612 VGND.t496 10.3303
R5739 VGND.n636 VGND.t245 10.3303
R5740 VGND.n660 VGND.t242 10.3303
R5741 VGND.n684 VGND.t87 10.3303
R5742 VGND.t117 VGND.n1069 10.3303
R5743 VGND.n1020 VGND.n1019 8.89919
R5744 VGND.n1051 VGND.n1028 8.89919
R5745 VGND.n1041 VGND.n1036 8.89919
R5746 VGND.n1745 VGND.n332 8.89919
R5747 VGND.n990 VGND.t4 7.40866
R5748 VGND.n771 VGND.t491 6.73519
R5749 VGND.n1771 VGND 6.60769
R5750 VGND.n1747 VGND.n137 6.22424
R5751 VGND.n1748 VGND.n1747 6.06172
R5752 VGND.n1732 VGND.n513 5.90952
R5753 VGND.n515 VGND.t325 5.8005
R5754 VGND.n515 VGND.t327 5.8005
R5755 VGND.n1280 VGND.t453 5.8005
R5756 VGND.n1280 VGND.t230 5.8005
R5757 VGND.n1279 VGND.t443 5.8005
R5758 VGND.n1279 VGND.t160 5.8005
R5759 VGND.n1278 VGND.t199 5.8005
R5760 VGND.n1278 VGND.t444 5.8005
R5761 VGND.n1276 VGND.t144 5.8005
R5762 VGND.n1276 VGND.t445 5.8005
R5763 VGND.n1275 VGND.t456 5.8005
R5764 VGND.n1275 VGND.t198 5.8005
R5765 VGND.n1273 VGND.t326 5.8005
R5766 VGND.n1273 VGND.t440 5.8005
R5767 VGND.n1272 VGND.t235 5.8005
R5768 VGND.n1272 VGND.t513 5.8005
R5769 VGND.n1270 VGND.t229 5.8005
R5770 VGND.n1270 VGND.t490 5.8005
R5771 VGND.n1269 VGND.t436 5.8005
R5772 VGND.n1269 VGND.t439 5.8005
R5773 VGND.n1224 VGND.t442 5.8005
R5774 VGND.n1224 VGND.t338 5.8005
R5775 VGND.n1225 VGND.t337 5.8005
R5776 VGND.n1225 VGND.t227 5.8005
R5777 VGND.n1238 VGND.t161 5.8005
R5778 VGND.n1238 VGND.t441 5.8005
R5779 VGND.n1255 VGND.t446 5.8005
R5780 VGND.n1255 VGND.t485 5.8005
R5781 VGND.n569 VGND.t512 5.8005
R5782 VGND.n569 VGND.t236 5.8005
R5783 VGND.n568 VGND.t438 5.8005
R5784 VGND.n568 VGND.t547 5.8005
R5785 VGND.n582 VGND.n564 5.54333
R5786 VGND.n1129 VGND.n592 5.54333
R5787 VGND.n608 VGND.n607 5.54333
R5788 VGND.n1116 VGND.n616 5.54333
R5789 VGND.n632 VGND.n631 5.54333
R5790 VGND.n1103 VGND.n640 5.54333
R5791 VGND.n656 VGND.n655 5.54333
R5792 VGND.n1090 VGND.n664 5.54333
R5793 VGND.n680 VGND.n679 5.54333
R5794 VGND.n1077 VGND.n688 5.54333
R5795 VGND.n1070 VGND.n698 5.54333
R5796 VGND.n725 VGND.n715 5.54333
R5797 VGND.t76 VGND.n1168 5.45827
R5798 VGND.n990 VGND.t124 5.16377
R5799 VGND VGND.n1771 4.64147
R5800 VGND.n1769 VGND.n1768 4.6393
R5801 VGND.n1139 VGND.n1138 3.89165
R5802 VGND.n1732 VGND.n1731 3.78262
R5803 VGND.t0 VGND.n137 3.70013
R5804 VGND VGND.n1802 3.50128
R5805 VGND.n295 VGND.n285 3.46248
R5806 VGND.n299 VGND.n298 3.46248
R5807 VGND.n291 VGND.n290 3.46248
R5808 VGND.n294 VGND.n286 3.46248
R5809 VGND.n276 VGND.n212 3.46248
R5810 VGND.n280 VGND.n279 3.46248
R5811 VGND.n272 VGND.n271 3.46248
R5812 VGND.n275 VGND.n213 3.46248
R5813 VGND.n243 VGND.n0 3.46248
R5814 VGND.n246 VGND.n235 3.46248
R5815 VGND.n149 VGND.n148 3.46248
R5816 VGND.n992 VGND.n741 3.46248
R5817 VGND.n995 VGND.n738 3.46248
R5818 VGND.n983 VGND.n765 3.46248
R5819 VGND.n987 VGND.n986 3.46248
R5820 VGND.n965 VGND.n964 3.46248
R5821 VGND.n968 VGND.n795 3.46248
R5822 VGND.n960 VGND.n959 3.46248
R5823 VGND.n963 VGND.n798 3.46248
R5824 VGND.n943 VGND.n942 3.46248
R5825 VGND.n946 VGND.n809 3.46248
R5826 VGND.n938 VGND.n937 3.46248
R5827 VGND.n941 VGND.n812 3.46248
R5828 VGND.n921 VGND.n920 3.46248
R5829 VGND.n924 VGND.n823 3.46248
R5830 VGND.n916 VGND.n915 3.46248
R5831 VGND.n919 VGND.n826 3.46248
R5832 VGND.n899 VGND.n898 3.46248
R5833 VGND.n902 VGND.n837 3.46248
R5834 VGND.n894 VGND.n893 3.46248
R5835 VGND.n897 VGND.n840 3.46248
R5836 VGND.n877 VGND.n876 3.46248
R5837 VGND.n880 VGND.n851 3.46248
R5838 VGND.n872 VGND.n871 3.46248
R5839 VGND.n875 VGND.n854 3.46248
R5840 VGND.n1774 VGND.n1772 3.46248
R5841 VGND.n127 VGND.n125 3.46248
R5842 VGND.n121 VGND.n119 3.46248
R5843 VGND.n115 VGND.n113 3.46248
R5844 VGND.n109 VGND.n107 3.46248
R5845 VGND.n103 VGND.n101 3.46248
R5846 VGND.n97 VGND.n95 3.46248
R5847 VGND.n91 VGND.n89 3.46248
R5848 VGND.n86 VGND.n68 3.46248
R5849 VGND.n1805 VGND.n1803 3.46248
R5850 VGND.n65 VGND.n63 3.46248
R5851 VGND.n59 VGND.n57 3.46248
R5852 VGND.n53 VGND.n51 3.46248
R5853 VGND.n47 VGND.n45 3.46248
R5854 VGND.n41 VGND.n39 3.46248
R5855 VGND.n35 VGND.n33 3.46248
R5856 VGND.n29 VGND.n27 3.46248
R5857 VGND.n23 VGND.n21 3.46248
R5858 VGND.n472 VGND.n471 3.46248
R5859 VGND.n469 VGND.n467 3.46248
R5860 VGND.n463 VGND.n461 3.46248
R5861 VGND.n457 VGND.n455 3.46248
R5862 VGND.n451 VGND.n449 3.46248
R5863 VGND.n445 VGND.n443 3.46248
R5864 VGND.n439 VGND.n437 3.46248
R5865 VGND.n433 VGND.n431 3.46248
R5866 VGND.n427 VGND.n425 3.46248
R5867 VGND.n421 VGND.n419 3.46248
R5868 VGND.n415 VGND.n413 3.46248
R5869 VGND.n409 VGND.n407 3.46248
R5870 VGND.n403 VGND.n401 3.46248
R5871 VGND.n397 VGND.n395 3.46248
R5872 VGND.n391 VGND.n389 3.46248
R5873 VGND.n385 VGND.n383 3.46248
R5874 VGND.n379 VGND.n377 3.46248
R5875 VGND.n374 VGND.n367 3.46248
R5876 VGND.n370 VGND.n369 3.46248
R5877 VGND.n513 VGND.n340 3.46248
R5878 VGND.n154 VGND.n153 3.46248
R5879 VGND.n1769 VGND.n4 3.07882
R5880 VGND.n1770 VGND.n1769 3.02279
R5881 VGND.n1706 VGND.n1705 3.0154
R5882 VGND.n1731 VGND 2.95362
R5883 VGND.n1750 VGND.n164 2.913
R5884 VGND.n1758 VGND.n1757 2.913
R5885 VGND.n257 VGND.n221 2.913
R5886 VGND.n253 VGND.n229 2.913
R5887 VGND.n323 VGND.n175 2.82278
R5888 VGND.n319 VGND.n181 2.82278
R5889 VGND.n322 VGND.n176 2.82278
R5890 VGND.n309 VGND.n195 2.82278
R5891 VGND.n289 VGND.n194 2.82278
R5892 VGND.n305 VGND.n203 2.82278
R5893 VGND.n308 VGND.n199 2.82278
R5894 VGND.n1011 VGND.n732 2.82278
R5895 VGND.n1007 VGND.n996 2.82278
R5896 VGND.n1010 VGND.n733 2.82278
R5897 VGND.n978 VGND.n769 2.82278
R5898 VGND.n982 VGND.n766 2.82278
R5899 VGND.n969 VGND.n794 2.82278
R5900 VGND.n973 VGND.n972 2.82278
R5901 VGND.n954 VGND.n952 2.82278
R5902 VGND.n958 VGND.n801 2.82278
R5903 VGND.n948 VGND.n947 2.82278
R5904 VGND.n951 VGND.n804 2.82278
R5905 VGND.n932 VGND.n930 2.82278
R5906 VGND.n936 VGND.n815 2.82278
R5907 VGND.n926 VGND.n925 2.82278
R5908 VGND.n929 VGND.n818 2.82278
R5909 VGND.n910 VGND.n908 2.82278
R5910 VGND.n914 VGND.n829 2.82278
R5911 VGND.n904 VGND.n903 2.82278
R5912 VGND.n907 VGND.n832 2.82278
R5913 VGND.n888 VGND.n886 2.82278
R5914 VGND.n892 VGND.n843 2.82278
R5915 VGND.n882 VGND.n881 2.82278
R5916 VGND.n885 VGND.n846 2.82278
R5917 VGND.n1015 VGND.n1014 2.82278
R5918 VGND.n327 VGND.n326 2.82278
R5919 VGND.n1801 VGND.n69 2.768
R5920 VGND.n1644 VGND.n74 2.768
R5921 VGND.n1658 VGND.n1645 2.768
R5922 VGND.n1663 VGND.n1634 2.768
R5923 VGND.n1664 VGND.n1633 2.768
R5924 VGND.n1671 VGND.n1670 2.768
R5925 VGND.n1676 VGND.n1618 2.768
R5926 VGND.n1681 VGND.n1610 2.768
R5927 VGND.n1682 VGND.n1609 2.768
R5928 VGND.n1689 VGND.n1688 2.768
R5929 VGND.n1694 VGND.n1594 2.768
R5930 VGND.n1699 VGND.n1586 2.768
R5931 VGND.n1700 VGND.n1585 2.768
R5932 VGND.n1531 VGND.n1530 2.768
R5933 VGND.n1542 VGND.n1523 2.768
R5934 VGND.n1544 VGND.n1543 2.768
R5935 VGND.n1517 VGND.n1411 2.768
R5936 VGND.n1516 VGND.n1412 2.768
R5937 VGND.n1511 VGND.n1510 2.768
R5938 VGND.n1507 VGND.n1424 2.768
R5939 VGND.n1502 VGND.n1501 2.768
R5940 VGND.n1498 VGND.n1436 2.768
R5941 VGND.n1493 VGND.n1492 2.768
R5942 VGND.n1489 VGND.n1448 2.768
R5943 VGND.n1484 VGND.n1483 2.768
R5944 VGND.n1480 VGND.n1460 2.768
R5945 VGND.n1475 VGND.n1474 2.768
R5946 VGND.n1552 VGND.n1158 2.768
R5947 VGND.n1557 VGND.n1150 2.768
R5948 VGND.n1558 VGND.n1149 2.768
R5949 VGND.n1565 VGND.n1564 2.768
R5950 VGND.n1407 VGND.n1401 2.52995
R5951 VGND.n1418 VGND.n1417 2.52995
R5952 VGND.n1430 VGND.n1429 2.52995
R5953 VGND.n1442 VGND.n1441 2.52995
R5954 VGND.n1454 VGND.n1453 2.52995
R5955 VGND.n1466 VGND.n1465 2.52995
R5956 VGND.n1159 VGND.n1155 2.52995
R5957 VGND.n1145 VGND.n566 2.52995
R5958 VGND.n1646 VGND.n1639 2.52995
R5959 VGND.n1647 VGND.n1627 2.52995
R5960 VGND.n1619 VGND.n1615 2.52995
R5961 VGND.n1620 VGND.n1603 2.52995
R5962 VGND.n1595 VGND.n1591 2.52995
R5963 VGND.n1596 VGND.n1579 2.52995
R5964 VGND.n1537 VGND.n1533 2.52995
R5965 VGND.n1796 VGND.n75 2.52995
R5966 VGND.n1731 VGND 2.40675
R5967 VGND.n1140 VGND.n1139 2.3961
R5968 VGND.n1752 VGND.n164 2.3255
R5969 VGND.n1757 VGND.n1756 2.3255
R5970 VGND.n1775 VGND.n128 2.3255
R5971 VGND.n1777 VGND.n122 2.3255
R5972 VGND.n1779 VGND.n116 2.3255
R5973 VGND.n1781 VGND.n110 2.3255
R5974 VGND.n1783 VGND.n104 2.3255
R5975 VGND.n1785 VGND.n98 2.3255
R5976 VGND.n1787 VGND.n92 2.3255
R5977 VGND.n1789 VGND.n87 2.3255
R5978 VGND.n1806 VGND.n66 2.3255
R5979 VGND.n1808 VGND.n60 2.3255
R5980 VGND.n1810 VGND.n54 2.3255
R5981 VGND.n1812 VGND.n48 2.3255
R5982 VGND.n1814 VGND.n42 2.3255
R5983 VGND.n1816 VGND.n36 2.3255
R5984 VGND.n1818 VGND.n30 2.3255
R5985 VGND.n1820 VGND.n24 2.3255
R5986 VGND.n1822 VGND.n19 2.3255
R5987 VGND.n475 VGND.n474 2.3255
R5988 VGND.n477 VGND.n464 2.3255
R5989 VGND.n479 VGND.n458 2.3255
R5990 VGND.n481 VGND.n452 2.3255
R5991 VGND.n483 VGND.n446 2.3255
R5992 VGND.n485 VGND.n440 2.3255
R5993 VGND.n487 VGND.n434 2.3255
R5994 VGND.n489 VGND.n428 2.3255
R5995 VGND.n491 VGND.n422 2.3255
R5996 VGND.n493 VGND.n416 2.3255
R5997 VGND.n495 VGND.n410 2.3255
R5998 VGND.n497 VGND.n404 2.3255
R5999 VGND.n499 VGND.n398 2.3255
R6000 VGND.n501 VGND.n392 2.3255
R6001 VGND.n503 VGND.n386 2.3255
R6002 VGND.n505 VGND.n380 2.3255
R6003 VGND.n507 VGND.n375 2.3255
R6004 VGND.n372 VGND.n371 2.3255
R6005 VGND.n512 VGND.n511 2.3255
R6006 VGND.n265 VGND.n221 2.3255
R6007 VGND.n231 VGND.n229 2.3255
R6008 VGND.n985 VGND.n764 2.3255
R6009 VGND.n994 VGND.n993 2.3255
R6010 VGND.n962 VGND.n961 2.3255
R6011 VGND.n967 VGND.n966 2.3255
R6012 VGND.n940 VGND.n939 2.3255
R6013 VGND.n945 VGND.n944 2.3255
R6014 VGND.n918 VGND.n917 2.3255
R6015 VGND.n923 VGND.n922 2.3255
R6016 VGND.n896 VGND.n895 2.3255
R6017 VGND.n901 VGND.n900 2.3255
R6018 VGND.n874 VGND.n873 2.3255
R6019 VGND.n879 VGND.n878 2.3255
R6020 VGND.n144 VGND.n143 2.3255
R6021 VGND.n293 VGND.n292 2.3255
R6022 VGND.n297 VGND.n284 2.3255
R6023 VGND.n274 VGND.n273 2.3255
R6024 VGND.n278 VGND.n211 2.3255
R6025 VGND.n245 VGND.n244 2.3255
R6026 VGND.n1139 VGND.n573 2.28621
R6027 VGND.n239 VGND.n238 2.17513
R6028 VGND.n1832 VGND.n4 2.15467
R6029 VGND.n1768 VGND.n130 2.15467
R6030 VGND.n1835 VGND.n1 2.1305
R6031 VGND.n132 VGND.n131 2.1305
R6032 VGND.n1712 VGND.n537 2.07965
R6033 VGND.n869 VGND.n858 1.95084
R6034 VGND.n865 VGND.n141 1.95084
R6035 VGND.n269 VGND.n216 1.95084
R6036 VGND.n251 VGND.n250 1.95084
R6037 VGND.n1766 VGND.n1765 1.8605
R6038 VGND.n1834 VGND.n1833 1.8605
R6039 VGND.n1730 VGND.n514 1.56378
R6040 VGND.n1302 VGND.n1284 1.56378
R6041 VGND.n1327 VGND.n1309 1.56378
R6042 VGND.n1352 VGND.n1334 1.56378
R6043 VGND.n1377 VGND.n1359 1.56378
R6044 VGND.n1387 VGND.n1384 1.56378
R6045 VGND.n1262 VGND.n1237 1.56378
R6046 VGND.n1723 VGND.n532 1.56378
R6047 VGND.n270 VGND.n269 1.52133
R6048 VGND VGND.n1557 1.3768
R6049 VGND.n1474 VGND 1.3768
R6050 VGND.n1483 VGND 1.3768
R6051 VGND.n1492 VGND 1.3768
R6052 VGND.n1501 VGND 1.3768
R6053 VGND.n1510 VGND 1.3768
R6054 VGND.n1517 VGND 1.3768
R6055 VGND VGND.n1542 1.3768
R6056 VGND.n1283 VGND.n517 1.37182
R6057 VGND.n1308 VGND.n1277 1.37182
R6058 VGND.n1333 VGND.n1274 1.37182
R6059 VGND.n1358 VGND.n1271 1.37182
R6060 VGND.n1383 VGND.n1268 1.37182
R6061 VGND.n1263 VGND.n1234 1.37182
R6062 VGND.n1259 VGND.n1258 1.37182
R6063 VGND.n573 VGND.n530 1.37182
R6064 VGND.n1009 VGND.n1008 1.32907
R6065 VGND.n1012 VGND.n727 1.32907
R6066 VGND.n971 VGND.n791 1.32907
R6067 VGND.n980 VGND.n979 1.32907
R6068 VGND.n950 VGND.n949 1.32907
R6069 VGND.n956 VGND.n955 1.32907
R6070 VGND.n928 VGND.n927 1.32907
R6071 VGND.n934 VGND.n933 1.32907
R6072 VGND.n906 VGND.n905 1.32907
R6073 VGND.n912 VGND.n911 1.32907
R6074 VGND.n884 VGND.n883 1.32907
R6075 VGND.n890 VGND.n889 1.32907
R6076 VGND.n321 VGND.n320 1.32907
R6077 VGND.n324 VGND.n170 1.32907
R6078 VGND.n307 VGND.n306 1.32907
R6079 VGND.n311 VGND.n310 1.32907
R6080 VGND.n870 VGND.n869 1.30085
R6081 VGND.n1140 VGND 1.21891
R6082 VGND.n1014 VGND.n729 0.959726
R6083 VGND.n326 VGND.n172 0.959726
R6084 VGND.n249 VGND.n234 0.957022
R6085 VGND.n268 VGND.n218 0.957022
R6086 VGND.n864 VGND.n862 0.957022
R6087 VGND.n868 VGND.n860 0.957022
R6088 VGND.n532 VGND.n531 0.785098
R6089 VGND.n1262 VGND.n1261 0.785098
R6090 VGND.n1384 VGND.n1267 0.785098
R6091 VGND.n1379 VGND.n1359 0.785098
R6092 VGND.n1354 VGND.n1334 0.785098
R6093 VGND.n1329 VGND.n1309 0.785098
R6094 VGND.n1304 VGND.n1284 0.785098
R6095 VGND.n1730 VGND.n1729 0.785098
R6096 VGND.n1771 VGND.n1770 0.738047
R6097 VGND.n202 VGND.n201 0.685283
R6098 VGND.n198 VGND.n197 0.685283
R6099 VGND.n179 VGND.n178 0.685283
R6100 VGND.n325 VGND.n174 0.685283
R6101 VGND.n849 VGND.n848 0.685283
R6102 VGND.n891 VGND.n845 0.685283
R6103 VGND.n835 VGND.n834 0.685283
R6104 VGND.n913 VGND.n831 0.685283
R6105 VGND.n821 VGND.n820 0.685283
R6106 VGND.n935 VGND.n817 0.685283
R6107 VGND.n807 VGND.n806 0.685283
R6108 VGND.n957 VGND.n803 0.685283
R6109 VGND.n970 VGND.n793 0.685283
R6110 VGND.n981 VGND.n768 0.685283
R6111 VGND.n736 VGND.n735 0.685283
R6112 VGND.n1013 VGND.n731 0.685283
R6113 VGND VGND.n1125 0.669618
R6114 VGND VGND.n1112 0.669618
R6115 VGND VGND.n1099 0.669618
R6116 VGND VGND.n1086 0.669618
R6117 VGND VGND.n1073 0.669618
R6118 VGND VGND.n1060 0.669618
R6119 VGND VGND.n1047 0.669618
R6120 VGND.n1798 VGND.n1797 0.58175
R6121 VGND.n1660 VGND.n1659 0.58175
R6122 VGND.n1667 VGND.n1628 0.58175
R6123 VGND.n1678 VGND.n1677 0.58175
R6124 VGND.n1685 VGND.n1604 0.58175
R6125 VGND.n1696 VGND.n1695 0.58175
R6126 VGND.n1703 VGND.n1580 0.58175
R6127 VGND.n1539 VGND.n1538 0.58175
R6128 VGND.n1520 VGND.n1402 0.58175
R6129 VGND.n1513 VGND.n1512 0.58175
R6130 VGND.n1504 VGND.n1503 0.58175
R6131 VGND.n1495 VGND.n1494 0.58175
R6132 VGND.n1486 VGND.n1485 0.58175
R6133 VGND.n1477 VGND.n1476 0.58175
R6134 VGND.n1554 VGND.n1553 0.58175
R6135 VGND.n1561 VGND.n567 0.58175
R6136 VGND.n1037 VGND.n338 0.58175
R6137 VGND.n1057 VGND.n1056 0.58175
R6138 VGND.n1083 VGND.n1082 0.58175
R6139 VGND.n1096 VGND.n1095 0.58175
R6140 VGND.n1109 VGND.n1108 0.58175
R6141 VGND.n1122 VGND.n1121 0.58175
R6142 VGND.n1135 VGND.n1134 0.58175
R6143 VGND.n1066 VGND.n1065 0.58175
R6144 VGND.n729 VGND 0.578086
R6145 VGND.n172 VGND 0.578086
R6146 VGND.n1564 VGND.n1140 0.53826
R6147 VGND VGND.n154 0.523938
R6148 VGND VGND.n246 0.523938
R6149 VGND VGND.n532 0.522821
R6150 VGND VGND.n1262 0.522821
R6151 VGND.n1384 VGND 0.522821
R6152 VGND.n1359 VGND 0.522821
R6153 VGND.n1334 VGND 0.522821
R6154 VGND.n1309 VGND 0.522821
R6155 VGND.n1284 VGND 0.522821
R6156 VGND VGND.n1730 0.522821
R6157 VGND.n1729 VGND.n1728 0.517167
R6158 VGND.n1304 VGND.n1303 0.517167
R6159 VGND.n1329 VGND.n1328 0.517167
R6160 VGND.n1354 VGND.n1353 0.517167
R6161 VGND.n1379 VGND.n1378 0.517167
R6162 VGND.n1267 VGND.n1223 0.517167
R6163 VGND.n1261 VGND.n1260 0.517167
R6164 VGND.n1724 VGND.n531 0.517167
R6165 VGND.n983 VGND 0.479667
R6166 VGND.n959 VGND 0.479667
R6167 VGND.n937 VGND 0.479667
R6168 VGND.n915 VGND 0.479667
R6169 VGND.n893 VGND 0.479667
R6170 VGND.n290 VGND 0.479667
R6171 VGND VGND.n995 0.466646
R6172 VGND VGND.n968 0.466646
R6173 VGND VGND.n946 0.466646
R6174 VGND VGND.n924 0.466646
R6175 VGND VGND.n902 0.466646
R6176 VGND VGND.n880 0.466646
R6177 VGND.n298 VGND 0.466646
R6178 VGND.n279 VGND 0.466646
R6179 VGND.n148 VGND 0.463123
R6180 VGND VGND.n0 0.463123
R6181 VGND.n1258 VGND 0.455857
R6182 VGND.n1263 VGND 0.455857
R6183 VGND VGND.n1383 0.455857
R6184 VGND VGND.n1358 0.455857
R6185 VGND VGND.n1333 0.455857
R6186 VGND VGND.n1308 0.455857
R6187 VGND VGND.n1283 0.455857
R6188 VGND.n866 VGND.n164 0.440404
R6189 VGND.n1757 VGND.n155 0.440404
R6190 VGND.n221 VGND.n219 0.440404
R6191 VGND.n247 VGND.n229 0.440404
R6192 VGND.n1011 VGND.n1010 0.430188
R6193 VGND.n972 VGND.n769 0.430188
R6194 VGND.n952 VGND.n951 0.430188
R6195 VGND.n930 VGND.n929 0.430188
R6196 VGND.n908 VGND.n907 0.430188
R6197 VGND.n886 VGND.n885 0.430188
R6198 VGND.n323 VGND.n322 0.430188
R6199 VGND.n309 VGND.n308 0.430188
R6200 VGND.n1802 VGND 0.426281
R6201 VGND.n863 VGND.n156 0.423227
R6202 VGND.n867 VGND.n163 0.423227
R6203 VGND.n248 VGND.n232 0.423227
R6204 VGND.n267 VGND.n266 0.423227
R6205 VGND.n271 VGND.n270 0.383313
R6206 VGND.n1037 VGND.n336 0.376971
R6207 VGND.n1056 VGND.n1055 0.376971
R6208 VGND.n1082 VGND.n1081 0.376971
R6209 VGND.n1095 VGND.n1094 0.376971
R6210 VGND.n1108 VGND.n1107 0.376971
R6211 VGND.n1121 VGND.n1120 0.376971
R6212 VGND.n1134 VGND.n1133 0.376971
R6213 VGND.n1066 VGND.n700 0.376971
R6214 VGND.n1012 VGND.n1011 0.359875
R6215 VGND.n1010 VGND.n1009 0.359875
R6216 VGND.n980 VGND.n769 0.359875
R6217 VGND.n972 VGND.n971 0.359875
R6218 VGND.n956 VGND.n952 0.359875
R6219 VGND.n951 VGND.n950 0.359875
R6220 VGND.n934 VGND.n930 0.359875
R6221 VGND.n929 VGND.n928 0.359875
R6222 VGND.n912 VGND.n908 0.359875
R6223 VGND.n907 VGND.n906 0.359875
R6224 VGND.n890 VGND.n886 0.359875
R6225 VGND.n885 VGND.n884 0.359875
R6226 VGND.n324 VGND.n323 0.359875
R6227 VGND.n322 VGND.n321 0.359875
R6228 VGND.n310 VGND.n309 0.359875
R6229 VGND.n308 VGND.n307 0.359875
R6230 VGND.n1137 VGND.n1136 0.324029
R6231 VGND.n595 VGND.n594 0.324029
R6232 VGND.n1124 VGND.n1123 0.324029
R6233 VGND.n619 VGND.n618 0.324029
R6234 VGND.n1111 VGND.n1110 0.324029
R6235 VGND.n643 VGND.n642 0.324029
R6236 VGND.n1098 VGND.n1097 0.324029
R6237 VGND.n667 VGND.n666 0.324029
R6238 VGND.n1085 VGND.n1084 0.324029
R6239 VGND.n691 VGND.n690 0.324029
R6240 VGND.n701 VGND.n693 0.324029
R6241 VGND.n1063 VGND.n1062 0.324029
R6242 VGND.n1059 VGND.n1058 0.324029
R6243 VGND.n1031 VGND.n1030 0.324029
R6244 VGND.n1046 VGND.n1045 0.324029
R6245 VGND.n1735 VGND.n1734 0.324029
R6246 VGND.n871 VGND.n870 0.323417
R6247 VGND.n866 VGND 0.306056
R6248 VGND.n155 VGND 0.306056
R6249 VGND VGND.n219 0.306056
R6250 VGND.n247 VGND 0.306056
R6251 VGND.n1770 VGND 0.284263
R6252 VGND.n1704 VGND.n1703 0.247896
R6253 VGND.n1703 VGND.n1702 0.247896
R6254 VGND.n1701 VGND.n1700 0.247896
R6255 VGND.n1699 VGND.n1698 0.247896
R6256 VGND.n1697 VGND.n1696 0.247896
R6257 VGND.n1696 VGND.n1590 0.247896
R6258 VGND.n1594 VGND.n1593 0.247896
R6259 VGND.n1688 VGND.n1687 0.247896
R6260 VGND.n1686 VGND.n1685 0.247896
R6261 VGND.n1685 VGND.n1684 0.247896
R6262 VGND.n1683 VGND.n1682 0.247896
R6263 VGND.n1681 VGND.n1680 0.247896
R6264 VGND.n1679 VGND.n1678 0.247896
R6265 VGND.n1678 VGND.n1614 0.247896
R6266 VGND.n1618 VGND.n1617 0.247896
R6267 VGND.n1670 VGND.n1669 0.247896
R6268 VGND.n1668 VGND.n1667 0.247896
R6269 VGND.n1667 VGND.n1666 0.247896
R6270 VGND.n1665 VGND.n1664 0.247896
R6271 VGND.n1663 VGND.n1662 0.247896
R6272 VGND.n1661 VGND.n1660 0.247896
R6273 VGND.n1660 VGND.n1638 0.247896
R6274 VGND.n1645 VGND.n1641 0.247896
R6275 VGND.n1644 VGND.n1643 0.247896
R6276 VGND.n1798 VGND.n73 0.247896
R6277 VGND.n1799 VGND.n1798 0.247896
R6278 VGND.n1801 VGND.n1800 0.247896
R6279 VGND.n1564 VGND.n1563 0.247896
R6280 VGND.n1562 VGND.n1561 0.247896
R6281 VGND.n1561 VGND.n1560 0.247896
R6282 VGND.n1559 VGND.n1558 0.247896
R6283 VGND.n1557 VGND.n1556 0.247896
R6284 VGND.n1555 VGND.n1554 0.247896
R6285 VGND.n1554 VGND.n1154 0.247896
R6286 VGND.n1158 VGND.n1157 0.247896
R6287 VGND.n1474 VGND.n1473 0.247896
R6288 VGND.n1477 VGND.n1464 0.247896
R6289 VGND.n1478 VGND.n1477 0.247896
R6290 VGND.n1480 VGND.n1479 0.247896
R6291 VGND.n1483 VGND.n1482 0.247896
R6292 VGND.n1486 VGND.n1452 0.247896
R6293 VGND.n1487 VGND.n1486 0.247896
R6294 VGND.n1489 VGND.n1488 0.247896
R6295 VGND.n1492 VGND.n1491 0.247896
R6296 VGND.n1495 VGND.n1440 0.247896
R6297 VGND.n1496 VGND.n1495 0.247896
R6298 VGND.n1498 VGND.n1497 0.247896
R6299 VGND.n1501 VGND.n1500 0.247896
R6300 VGND.n1504 VGND.n1428 0.247896
R6301 VGND.n1505 VGND.n1504 0.247896
R6302 VGND.n1507 VGND.n1506 0.247896
R6303 VGND.n1510 VGND.n1509 0.247896
R6304 VGND.n1513 VGND.n1416 0.247896
R6305 VGND.n1514 VGND.n1513 0.247896
R6306 VGND.n1516 VGND.n1515 0.247896
R6307 VGND.n1518 VGND.n1517 0.247896
R6308 VGND.n1520 VGND.n1519 0.247896
R6309 VGND.n1521 VGND.n1520 0.247896
R6310 VGND.n1543 VGND.n1522 0.247896
R6311 VGND.n1542 VGND.n1541 0.247896
R6312 VGND.n1540 VGND.n1539 0.247896
R6313 VGND.n1539 VGND.n1527 0.247896
R6314 VGND.n1530 VGND.n1529 0.247896
R6315 VGND.n570 VGND.n531 0.246036
R6316 VGND.n1261 VGND.n1239 0.246036
R6317 VGND.n1267 VGND.n1266 0.246036
R6318 VGND.n1380 VGND.n1379 0.246036
R6319 VGND.n1355 VGND.n1354 0.246036
R6320 VGND.n1330 VGND.n1329 0.246036
R6321 VGND.n1305 VGND.n1304 0.246036
R6322 VGND.n1729 VGND.n516 0.246036
R6323 VGND.n1138 VGND.n1137 0.239471
R6324 VGND.n1125 VGND.n1124 0.239471
R6325 VGND.n1112 VGND.n1111 0.239471
R6326 VGND.n1099 VGND.n1098 0.239471
R6327 VGND.n1086 VGND.n1085 0.239471
R6328 VGND.n1073 VGND.n693 0.239471
R6329 VGND.n1060 VGND.n1059 0.239471
R6330 VGND.n1047 VGND.n1046 0.239471
R6331 VGND.n1126 VGND.n595 0.232118
R6332 VGND.n1113 VGND.n619 0.232118
R6333 VGND.n1100 VGND.n643 0.232118
R6334 VGND.n1087 VGND.n667 0.232118
R6335 VGND.n1074 VGND.n691 0.232118
R6336 VGND.n1062 VGND.n1061 0.232118
R6337 VGND.n1048 VGND.n1031 0.232118
R6338 VGND.n1734 VGND.n1733 0.232118
R6339 VGND.n1766 VGND.n131 0.230892
R6340 VGND.n1835 VGND.n1834 0.230892
R6341 VGND.n1705 VGND.n1704 0.229667
R6342 VGND.n1702 VGND.n1701 0.229667
R6343 VGND.n1698 VGND.n1697 0.229667
R6344 VGND.n1593 VGND.n1590 0.229667
R6345 VGND.n1687 VGND.n1686 0.229667
R6346 VGND.n1684 VGND.n1683 0.229667
R6347 VGND.n1680 VGND.n1679 0.229667
R6348 VGND.n1617 VGND.n1614 0.229667
R6349 VGND.n1669 VGND.n1668 0.229667
R6350 VGND.n1666 VGND.n1665 0.229667
R6351 VGND.n1662 VGND.n1661 0.229667
R6352 VGND.n1641 VGND.n1638 0.229667
R6353 VGND.n1643 VGND.n73 0.229667
R6354 VGND.n1800 VGND.n1799 0.229667
R6355 VGND.n1563 VGND.n1562 0.229667
R6356 VGND.n1560 VGND.n1559 0.229667
R6357 VGND.n1556 VGND.n1555 0.229667
R6358 VGND.n1157 VGND.n1154 0.229667
R6359 VGND.n1473 VGND.n1464 0.229667
R6360 VGND.n1479 VGND.n1478 0.229667
R6361 VGND.n1482 VGND.n1452 0.229667
R6362 VGND.n1488 VGND.n1487 0.229667
R6363 VGND.n1491 VGND.n1440 0.229667
R6364 VGND.n1497 VGND.n1496 0.229667
R6365 VGND.n1500 VGND.n1428 0.229667
R6366 VGND.n1506 VGND.n1505 0.229667
R6367 VGND.n1509 VGND.n1416 0.229667
R6368 VGND.n1515 VGND.n1514 0.229667
R6369 VGND.n1519 VGND.n1518 0.229667
R6370 VGND.n1522 VGND.n1521 0.229667
R6371 VGND.n1541 VGND.n1540 0.229667
R6372 VGND.n1529 VGND.n1527 0.229667
R6373 VGND.n1013 VGND.n1012 0.229667
R6374 VGND.n1009 VGND.n736 0.229667
R6375 VGND.n981 VGND.n980 0.229667
R6376 VGND.n971 VGND.n970 0.229667
R6377 VGND.n957 VGND.n956 0.229667
R6378 VGND.n950 VGND.n807 0.229667
R6379 VGND.n935 VGND.n934 0.229667
R6380 VGND.n928 VGND.n821 0.229667
R6381 VGND.n913 VGND.n912 0.229667
R6382 VGND.n906 VGND.n835 0.229667
R6383 VGND.n891 VGND.n890 0.229667
R6384 VGND.n884 VGND.n849 0.229667
R6385 VGND.n325 VGND.n324 0.229667
R6386 VGND.n321 VGND.n179 0.229667
R6387 VGND.n310 VGND.n198 0.229667
R6388 VGND.n307 VGND.n202 0.229667
R6389 VGND.n781 VGND.t4 0.22499
R6390 VGND.n1802 VGND.n68 0.212219
R6391 VGND.n572 VGND.n571 0.196929
R6392 VGND.n571 VGND.n570 0.196929
R6393 VGND.n1257 VGND.n1256 0.196929
R6394 VGND.n1256 VGND.n1239 0.196929
R6395 VGND.n1265 VGND.n1264 0.196929
R6396 VGND.n1266 VGND.n1265 0.196929
R6397 VGND.n1382 VGND.n1381 0.196929
R6398 VGND.n1381 VGND.n1380 0.196929
R6399 VGND.n1357 VGND.n1356 0.196929
R6400 VGND.n1356 VGND.n1355 0.196929
R6401 VGND.n1332 VGND.n1331 0.196929
R6402 VGND.n1331 VGND.n1330 0.196929
R6403 VGND.n1307 VGND.n1306 0.196929
R6404 VGND.n1306 VGND.n1305 0.196929
R6405 VGND.n1282 VGND.n1281 0.196929
R6406 VGND.n1281 VGND.n516 0.196929
R6407 VGND VGND.n982 0.191906
R6408 VGND VGND.n958 0.191906
R6409 VGND VGND.n936 0.191906
R6410 VGND VGND.n914 0.191906
R6411 VGND VGND.n892 0.191906
R6412 VGND VGND.n289 0.191906
R6413 VGND.n87 VGND.n68 0.189302
R6414 VGND.n92 VGND.n91 0.189302
R6415 VGND.n98 VGND.n97 0.189302
R6416 VGND.n104 VGND.n103 0.189302
R6417 VGND.n110 VGND.n109 0.189302
R6418 VGND.n116 VGND.n115 0.189302
R6419 VGND.n122 VGND.n121 0.189302
R6420 VGND.n128 VGND.n127 0.189302
R6421 VGND.n513 VGND.n512 0.189302
R6422 VGND.n372 VGND.n370 0.189302
R6423 VGND.n375 VGND.n374 0.189302
R6424 VGND.n380 VGND.n379 0.189302
R6425 VGND.n386 VGND.n385 0.189302
R6426 VGND.n392 VGND.n391 0.189302
R6427 VGND.n398 VGND.n397 0.189302
R6428 VGND.n404 VGND.n403 0.189302
R6429 VGND.n410 VGND.n409 0.189302
R6430 VGND.n416 VGND.n415 0.189302
R6431 VGND.n422 VGND.n421 0.189302
R6432 VGND.n428 VGND.n427 0.189302
R6433 VGND.n434 VGND.n433 0.189302
R6434 VGND.n440 VGND.n439 0.189302
R6435 VGND.n446 VGND.n445 0.189302
R6436 VGND.n452 VGND.n451 0.189302
R6437 VGND.n458 VGND.n457 0.189302
R6438 VGND.n464 VGND.n463 0.189302
R6439 VGND.n474 VGND.n469 0.189302
R6440 VGND.n472 VGND.n19 0.189302
R6441 VGND.n24 VGND.n23 0.189302
R6442 VGND.n30 VGND.n29 0.189302
R6443 VGND.n36 VGND.n35 0.189302
R6444 VGND.n42 VGND.n41 0.189302
R6445 VGND.n48 VGND.n47 0.189302
R6446 VGND.n54 VGND.n53 0.189302
R6447 VGND.n60 VGND.n59 0.189302
R6448 VGND.n66 VGND.n65 0.189302
R6449 VGND.n995 VGND.n994 0.189302
R6450 VGND.n986 VGND.n985 0.189302
R6451 VGND.n968 VGND.n967 0.189302
R6452 VGND.n963 VGND.n962 0.189302
R6453 VGND.n946 VGND.n945 0.189302
R6454 VGND.n941 VGND.n940 0.189302
R6455 VGND.n924 VGND.n923 0.189302
R6456 VGND.n919 VGND.n918 0.189302
R6457 VGND.n902 VGND.n901 0.189302
R6458 VGND.n897 VGND.n896 0.189302
R6459 VGND.n880 VGND.n879 0.189302
R6460 VGND.n875 VGND.n874 0.189302
R6461 VGND.n154 VGND.n143 0.189302
R6462 VGND.n298 VGND.n297 0.189302
R6463 VGND.n294 VGND.n293 0.189302
R6464 VGND.n279 VGND.n278 0.189302
R6465 VGND.n275 VGND.n274 0.189302
R6466 VGND.n246 VGND.n245 0.189302
R6467 VGND VGND.n1732 0.172069
R6468 VGND.n869 VGND.n868 0.169771
R6469 VGND.n865 VGND.n864 0.169771
R6470 VGND.n269 VGND.n268 0.169771
R6471 VGND.n250 VGND.n249 0.169771
R6472 VGND.n868 VGND.n867 0.168035
R6473 VGND.n864 VGND.n863 0.168035
R6474 VGND.n268 VGND.n267 0.168035
R6475 VGND.n249 VGND.n248 0.168035
R6476 VGND VGND.n865 0.15675
R6477 VGND.n250 VGND 0.15675
R6478 VGND.n1700 VGND 0.147635
R6479 VGND VGND.n1594 0.147635
R6480 VGND.n1682 VGND 0.147635
R6481 VGND VGND.n1618 0.147635
R6482 VGND.n1664 VGND 0.147635
R6483 VGND.n1645 VGND 0.147635
R6484 VGND VGND.n1801 0.147635
R6485 VGND.n1558 VGND 0.147635
R6486 VGND VGND.n1158 0.147635
R6487 VGND VGND.n1480 0.147635
R6488 VGND VGND.n1489 0.147635
R6489 VGND VGND.n1498 0.147635
R6490 VGND VGND.n1507 0.147635
R6491 VGND VGND.n1516 0.147635
R6492 VGND.n1543 VGND 0.147635
R6493 VGND.n1530 VGND 0.147635
R6494 VGND.n573 VGND.n572 0.146705
R6495 VGND.n1258 VGND.n1257 0.146705
R6496 VGND.n1264 VGND.n1263 0.146705
R6497 VGND.n1383 VGND.n1382 0.146705
R6498 VGND.n1358 VGND.n1357 0.146705
R6499 VGND.n1333 VGND.n1332 0.146705
R6500 VGND.n1308 VGND.n1307 0.146705
R6501 VGND.n1283 VGND.n1282 0.146705
R6502 VGND.n986 VGND.n741 0.141125
R6503 VGND.n964 VGND.n963 0.141125
R6504 VGND.n942 VGND.n941 0.141125
R6505 VGND.n920 VGND.n919 0.141125
R6506 VGND.n898 VGND.n897 0.141125
R6507 VGND.n876 VGND.n875 0.141125
R6508 VGND.n295 VGND.n294 0.141125
R6509 VGND.n276 VGND.n275 0.141125
R6510 VGND.n91 VGND.n90 0.13201
R6511 VGND.n97 VGND.n96 0.13201
R6512 VGND.n103 VGND.n102 0.13201
R6513 VGND.n109 VGND.n108 0.13201
R6514 VGND.n115 VGND.n114 0.13201
R6515 VGND.n121 VGND.n120 0.13201
R6516 VGND.n127 VGND.n126 0.13201
R6517 VGND.n1772 VGND.n129 0.13201
R6518 VGND.n370 VGND.n341 0.13201
R6519 VGND.n374 VGND.n373 0.13201
R6520 VGND.n379 VGND.n378 0.13201
R6521 VGND.n385 VGND.n384 0.13201
R6522 VGND.n391 VGND.n390 0.13201
R6523 VGND.n397 VGND.n396 0.13201
R6524 VGND.n403 VGND.n402 0.13201
R6525 VGND.n409 VGND.n408 0.13201
R6526 VGND.n415 VGND.n414 0.13201
R6527 VGND.n421 VGND.n420 0.13201
R6528 VGND.n427 VGND.n426 0.13201
R6529 VGND.n433 VGND.n432 0.13201
R6530 VGND.n439 VGND.n438 0.13201
R6531 VGND.n445 VGND.n444 0.13201
R6532 VGND.n451 VGND.n450 0.13201
R6533 VGND.n457 VGND.n456 0.13201
R6534 VGND.n463 VGND.n462 0.13201
R6535 VGND.n469 VGND.n468 0.13201
R6536 VGND.n473 VGND.n472 0.13201
R6537 VGND.n23 VGND.n22 0.13201
R6538 VGND.n29 VGND.n28 0.13201
R6539 VGND.n35 VGND.n34 0.13201
R6540 VGND.n41 VGND.n40 0.13201
R6541 VGND.n47 VGND.n46 0.13201
R6542 VGND.n53 VGND.n52 0.13201
R6543 VGND.n59 VGND.n58 0.13201
R6544 VGND.n65 VGND.n64 0.13201
R6545 VGND.n1803 VGND.n67 0.13201
R6546 VGND.n741 VGND.n739 0.13201
R6547 VGND.n984 VGND.n983 0.13201
R6548 VGND.n964 VGND.n796 0.13201
R6549 VGND.n959 VGND.n799 0.13201
R6550 VGND.n942 VGND.n810 0.13201
R6551 VGND.n937 VGND.n813 0.13201
R6552 VGND.n920 VGND.n824 0.13201
R6553 VGND.n915 VGND.n827 0.13201
R6554 VGND.n898 VGND.n838 0.13201
R6555 VGND.n893 VGND.n841 0.13201
R6556 VGND.n876 VGND.n852 0.13201
R6557 VGND.n871 VGND.n855 0.13201
R6558 VGND.n148 VGND.n147 0.13201
R6559 VGND.n296 VGND.n295 0.13201
R6560 VGND.n290 VGND.n287 0.13201
R6561 VGND.n277 VGND.n276 0.13201
R6562 VGND.n271 VGND.n214 0.13201
R6563 VGND.n236 VGND.n0 0.13201
R6564 VGND.n996 VGND.n736 0.130708
R6565 VGND.n970 VGND.n969 0.130708
R6566 VGND.n947 VGND.n807 0.130708
R6567 VGND.n925 VGND.n821 0.130708
R6568 VGND.n903 VGND.n835 0.130708
R6569 VGND.n881 VGND.n849 0.130708
R6570 VGND.n181 VGND.n179 0.130708
R6571 VGND.n203 VGND.n202 0.130708
R6572 VGND.n594 VGND.n576 0.124275
R6573 VGND.n618 VGND.n598 0.124275
R6574 VGND.n642 VGND.n622 0.124275
R6575 VGND.n666 VGND.n646 0.124275
R6576 VGND.n690 VGND.n670 0.124275
R6577 VGND.n1064 VGND.n1063 0.124275
R6578 VGND.n1030 VGND.n707 0.124275
R6579 VGND.n1736 VGND.n1735 0.124275
R6580 VGND VGND.n1013 0.124198
R6581 VGND VGND.n981 0.124198
R6582 VGND VGND.n957 0.124198
R6583 VGND VGND.n935 0.124198
R6584 VGND VGND.n913 0.124198
R6585 VGND VGND.n891 0.124198
R6586 VGND VGND.n325 0.124198
R6587 VGND VGND.n198 0.124198
R6588 VGND.n1768 VGND.n1767 0.121824
R6589 VGND.n4 VGND.n2 0.121824
R6590 VGND.n1136 VGND.n1135 0.120598
R6591 VGND.n1123 VGND.n1122 0.120598
R6592 VGND.n1110 VGND.n1109 0.120598
R6593 VGND.n1097 VGND.n1096 0.120598
R6594 VGND.n1084 VGND.n1083 0.120598
R6595 VGND.n1065 VGND.n701 0.120598
R6596 VGND.n1058 VGND.n1057 0.120598
R6597 VGND.n1045 VGND.n338 0.120598
R6598 VGND.n1126 VGND 0.113245
R6599 VGND.n1113 VGND 0.113245
R6600 VGND.n1100 VGND 0.113245
R6601 VGND.n1087 VGND 0.113245
R6602 VGND.n1074 VGND 0.113245
R6603 VGND.n1061 VGND 0.113245
R6604 VGND.n1048 VGND 0.113245
R6605 VGND.n1733 VGND 0.113245
R6606 VGND.n1767 VGND.n1766 0.108343
R6607 VGND.n1834 VGND.n2 0.108343
R6608 VGND.n867 VGND.n866 0.104667
R6609 VGND.n863 VGND.n155 0.104667
R6610 VGND.n267 VGND.n219 0.104667
R6611 VGND.n248 VGND.n247 0.104667
R6612 VGND VGND.n1699 0.0721146
R6613 VGND.n1688 VGND 0.0721146
R6614 VGND VGND.n1681 0.0721146
R6615 VGND.n1670 VGND 0.0721146
R6616 VGND VGND.n1663 0.0721146
R6617 VGND VGND.n1644 0.0721146
R6618 VGND.n1772 VGND 0.0708125
R6619 VGND.n1803 VGND 0.0708125
R6620 VGND.n996 VGND 0.0695104
R6621 VGND.n969 VGND 0.0695104
R6622 VGND.n947 VGND 0.0695104
R6623 VGND.n925 VGND 0.0695104
R6624 VGND.n903 VGND 0.0695104
R6625 VGND.n881 VGND 0.0695104
R6626 VGND VGND.n181 0.0695104
R6627 VGND VGND.n203 0.0695104
R6628 VGND.n90 VGND.n87 0.0577917
R6629 VGND.n96 VGND.n92 0.0577917
R6630 VGND.n102 VGND.n98 0.0577917
R6631 VGND.n108 VGND.n104 0.0577917
R6632 VGND.n114 VGND.n110 0.0577917
R6633 VGND.n120 VGND.n116 0.0577917
R6634 VGND.n126 VGND.n122 0.0577917
R6635 VGND.n129 VGND.n128 0.0577917
R6636 VGND.n512 VGND.n341 0.0577917
R6637 VGND.n373 VGND.n372 0.0577917
R6638 VGND.n378 VGND.n375 0.0577917
R6639 VGND.n384 VGND.n380 0.0577917
R6640 VGND.n390 VGND.n386 0.0577917
R6641 VGND.n396 VGND.n392 0.0577917
R6642 VGND.n402 VGND.n398 0.0577917
R6643 VGND.n408 VGND.n404 0.0577917
R6644 VGND.n414 VGND.n410 0.0577917
R6645 VGND.n420 VGND.n416 0.0577917
R6646 VGND.n426 VGND.n422 0.0577917
R6647 VGND.n432 VGND.n428 0.0577917
R6648 VGND.n438 VGND.n434 0.0577917
R6649 VGND.n444 VGND.n440 0.0577917
R6650 VGND.n450 VGND.n446 0.0577917
R6651 VGND.n456 VGND.n452 0.0577917
R6652 VGND.n462 VGND.n458 0.0577917
R6653 VGND.n468 VGND.n464 0.0577917
R6654 VGND.n474 VGND.n473 0.0577917
R6655 VGND.n22 VGND.n19 0.0577917
R6656 VGND.n28 VGND.n24 0.0577917
R6657 VGND.n34 VGND.n30 0.0577917
R6658 VGND.n40 VGND.n36 0.0577917
R6659 VGND.n46 VGND.n42 0.0577917
R6660 VGND.n52 VGND.n48 0.0577917
R6661 VGND.n58 VGND.n54 0.0577917
R6662 VGND.n64 VGND.n60 0.0577917
R6663 VGND.n67 VGND.n66 0.0577917
R6664 VGND.n994 VGND.n739 0.0577917
R6665 VGND.n985 VGND.n984 0.0577917
R6666 VGND.n967 VGND.n796 0.0577917
R6667 VGND.n962 VGND.n799 0.0577917
R6668 VGND.n945 VGND.n810 0.0577917
R6669 VGND.n940 VGND.n813 0.0577917
R6670 VGND.n923 VGND.n824 0.0577917
R6671 VGND.n918 VGND.n827 0.0577917
R6672 VGND.n901 VGND.n838 0.0577917
R6673 VGND.n896 VGND.n841 0.0577917
R6674 VGND.n879 VGND.n852 0.0577917
R6675 VGND.n874 VGND.n855 0.0577917
R6676 VGND.n147 VGND.n143 0.0577917
R6677 VGND.n297 VGND.n296 0.0577917
R6678 VGND.n293 VGND.n287 0.0577917
R6679 VGND.n278 VGND.n277 0.0577917
R6680 VGND.n274 VGND.n214 0.0577917
R6681 VGND.n245 VGND.n236 0.0577917
R6682 VGND.n729 VGND 0.0522857
R6683 VGND.n172 VGND 0.0522857
R6684 VGND.n270 VGND 0.0213333
R6685 VGND VGND.n131 0.0164314
R6686 VGND VGND.n1835 0.0164314
R6687 VGND.n870 VGND 0.00918056
R6688 VGND.n270 VGND 0.00918056
R6689 VGND.n1014 VGND 0.00701042
R6690 VGND.n982 VGND 0.00701042
R6691 VGND.n958 VGND 0.00701042
R6692 VGND.n936 VGND 0.00701042
R6693 VGND.n914 VGND 0.00701042
R6694 VGND.n892 VGND 0.00701042
R6695 VGND.n326 VGND 0.00701042
R6696 VGND.n289 VGND 0.00701042
R6697 VGND.n1135 VGND.n576 0.00417647
R6698 VGND.n1122 VGND.n598 0.00417647
R6699 VGND.n1109 VGND.n622 0.00417647
R6700 VGND.n1096 VGND.n646 0.00417647
R6701 VGND.n1083 VGND.n670 0.00417647
R6702 VGND.n1065 VGND.n1064 0.00417647
R6703 VGND.n1057 VGND.n707 0.00417647
R6704 VGND.n1736 VGND.n338 0.00417647
R6705 a_9330_16954.n1 a_9330_16954.t9 543.053
R6706 a_9330_16954.n2 a_9330_16954.t29 543.053
R6707 a_9330_16954.n4 a_9330_16954.t16 543.053
R6708 a_9330_16954.n6 a_9330_16954.t35 543.053
R6709 a_9330_16954.n8 a_9330_16954.t23 543.053
R6710 a_9330_16954.n10 a_9330_16954.t25 543.053
R6711 a_9330_16954.n12 a_9330_16954.t11 543.053
R6712 a_9330_16954.n14 a_9330_16954.t31 543.053
R6713 a_9330_16954.n16 a_9330_16954.t19 543.053
R6714 a_9330_16954.n18 a_9330_16954.t37 543.053
R6715 a_9330_16954.n20 a_9330_16954.t18 543.053
R6716 a_9330_16954.n22 a_9330_16954.t36 543.053
R6717 a_9330_16954.n24 a_9330_16954.t24 543.053
R6718 a_9330_16954.n26 a_9330_16954.t10 543.053
R6719 a_9330_16954.n28 a_9330_16954.t30 543.053
R6720 a_9330_16954.n0 a_9330_16954.t17 543.053
R6721 a_9330_16954.n1 a_9330_16954.t38 221.72
R6722 a_9330_16954.n2 a_9330_16954.t26 221.72
R6723 a_9330_16954.n4 a_9330_16954.t12 221.72
R6724 a_9330_16954.n6 a_9330_16954.t32 221.72
R6725 a_9330_16954.n8 a_9330_16954.t20 221.72
R6726 a_9330_16954.n10 a_9330_16954.t22 221.72
R6727 a_9330_16954.n12 a_9330_16954.t8 221.72
R6728 a_9330_16954.n14 a_9330_16954.t28 221.72
R6729 a_9330_16954.n16 a_9330_16954.t15 221.72
R6730 a_9330_16954.n18 a_9330_16954.t34 221.72
R6731 a_9330_16954.n20 a_9330_16954.t14 221.72
R6732 a_9330_16954.n22 a_9330_16954.t33 221.72
R6733 a_9330_16954.n24 a_9330_16954.t21 221.72
R6734 a_9330_16954.n26 a_9330_16954.t39 221.72
R6735 a_9330_16954.n28 a_9330_16954.t27 221.72
R6736 a_9330_16954.n0 a_9330_16954.t13 221.72
R6737 a_9330_16954.n3 a_9330_16954.n1 218.32
R6738 a_9330_16954.n3 a_9330_16954.n2 217.734
R6739 a_9330_16954.n5 a_9330_16954.n4 217.734
R6740 a_9330_16954.n7 a_9330_16954.n6 217.734
R6741 a_9330_16954.n9 a_9330_16954.n8 217.734
R6742 a_9330_16954.n11 a_9330_16954.n10 217.734
R6743 a_9330_16954.n13 a_9330_16954.n12 217.734
R6744 a_9330_16954.n15 a_9330_16954.n14 217.734
R6745 a_9330_16954.n17 a_9330_16954.n16 217.734
R6746 a_9330_16954.n19 a_9330_16954.n18 217.734
R6747 a_9330_16954.n21 a_9330_16954.n20 217.734
R6748 a_9330_16954.n23 a_9330_16954.n22 217.734
R6749 a_9330_16954.n25 a_9330_16954.n24 217.734
R6750 a_9330_16954.n27 a_9330_16954.n26 217.734
R6751 a_9330_16954.n29 a_9330_16954.n28 217.734
R6752 a_9330_16954.n30 a_9330_16954.n0 213.234
R6753 a_9330_16954.n33 a_9330_16954.t6 85.2499
R6754 a_9330_16954.n35 a_9330_16954.t5 85.2499
R6755 a_9330_16954.t7 a_9330_16954.n37 85.2499
R6756 a_9330_16954.n31 a_9330_16954.t4 84.7173
R6757 a_9330_16954.n37 a_9330_16954.t3 83.7172
R6758 a_9330_16954.n32 a_9330_16954.t0 83.7172
R6759 a_9330_16954.n33 a_9330_16954.t2 83.7172
R6760 a_9330_16954.n35 a_9330_16954.t1 83.7172
R6761 a_9330_16954.n34 a_9330_16954.n32 5.16238
R6762 a_9330_16954.n36 a_9330_16954.n35 5.16238
R6763 a_9330_16954.n30 a_9330_16954.n29 5.08518
R6764 a_9330_16954.n34 a_9330_16954.n33 4.64452
R6765 a_9330_16954.n37 a_9330_16954.n36 4.64452
R6766 a_9330_16954.n5 a_9330_16954.n3 0.585177
R6767 a_9330_16954.n7 a_9330_16954.n5 0.585177
R6768 a_9330_16954.n9 a_9330_16954.n7 0.585177
R6769 a_9330_16954.n11 a_9330_16954.n9 0.585177
R6770 a_9330_16954.n13 a_9330_16954.n11 0.585177
R6771 a_9330_16954.n15 a_9330_16954.n13 0.585177
R6772 a_9330_16954.n17 a_9330_16954.n15 0.585177
R6773 a_9330_16954.n19 a_9330_16954.n17 0.585177
R6774 a_9330_16954.n21 a_9330_16954.n19 0.585177
R6775 a_9330_16954.n23 a_9330_16954.n21 0.585177
R6776 a_9330_16954.n25 a_9330_16954.n23 0.585177
R6777 a_9330_16954.n27 a_9330_16954.n25 0.585177
R6778 a_9330_16954.n29 a_9330_16954.n27 0.585177
R6779 a_9330_16954.n36 a_9330_16954.n34 0.518357
R6780 a_9330_16954.n32 a_9330_16954.n31 0.36463
R6781 a_9330_16954.n31 a_9330_16954.n30 0.226306
R6782 tdc_0.vernier_delay_line_0.stop_strong.n52 tdc_0.vernier_delay_line_0.stop_strong.t86 851.506
R6783 tdc_0.vernier_delay_line_0.stop_strong.n45 tdc_0.vernier_delay_line_0.stop_strong.t48 851.506
R6784 tdc_0.vernier_delay_line_0.stop_strong.n38 tdc_0.vernier_delay_line_0.stop_strong.t76 851.506
R6785 tdc_0.vernier_delay_line_0.stop_strong.n31 tdc_0.vernier_delay_line_0.stop_strong.t66 851.506
R6786 tdc_0.vernier_delay_line_0.stop_strong.n24 tdc_0.vernier_delay_line_0.stop_strong.t49 851.506
R6787 tdc_0.vernier_delay_line_0.stop_strong.n17 tdc_0.vernier_delay_line_0.stop_strong.t61 851.506
R6788 tdc_0.vernier_delay_line_0.stop_strong.n10 tdc_0.vernier_delay_line_0.stop_strong.t80 851.506
R6789 tdc_0.vernier_delay_line_0.stop_strong.n4 tdc_0.vernier_delay_line_0.stop_strong.t56 851.506
R6790 tdc_0.vernier_delay_line_0.stop_strong.n52 tdc_0.vernier_delay_line_0.stop_strong.t79 850.414
R6791 tdc_0.vernier_delay_line_0.stop_strong.n45 tdc_0.vernier_delay_line_0.stop_strong.t58 850.414
R6792 tdc_0.vernier_delay_line_0.stop_strong.n38 tdc_0.vernier_delay_line_0.stop_strong.t74 850.414
R6793 tdc_0.vernier_delay_line_0.stop_strong.n31 tdc_0.vernier_delay_line_0.stop_strong.t77 850.414
R6794 tdc_0.vernier_delay_line_0.stop_strong.n24 tdc_0.vernier_delay_line_0.stop_strong.t45 850.414
R6795 tdc_0.vernier_delay_line_0.stop_strong.n17 tdc_0.vernier_delay_line_0.stop_strong.t59 850.414
R6796 tdc_0.vernier_delay_line_0.stop_strong.n10 tdc_0.vernier_delay_line_0.stop_strong.t39 850.414
R6797 tdc_0.vernier_delay_line_0.stop_strong.n4 tdc_0.vernier_delay_line_0.stop_strong.t87 850.414
R6798 tdc_0.vernier_delay_line_0.stop_strong.n48 tdc_0.vernier_delay_line_0.stop_strong.t75 641.061
R6799 tdc_0.vernier_delay_line_0.stop_strong.n41 tdc_0.vernier_delay_line_0.stop_strong.t38 641.061
R6800 tdc_0.vernier_delay_line_0.stop_strong.n34 tdc_0.vernier_delay_line_0.stop_strong.t81 641.061
R6801 tdc_0.vernier_delay_line_0.stop_strong.n27 tdc_0.vernier_delay_line_0.stop_strong.t70 641.061
R6802 tdc_0.vernier_delay_line_0.stop_strong.n20 tdc_0.vernier_delay_line_0.stop_strong.t40 641.061
R6803 tdc_0.vernier_delay_line_0.stop_strong.n13 tdc_0.vernier_delay_line_0.stop_strong.t52 641.061
R6804 tdc_0.vernier_delay_line_0.stop_strong.n6 tdc_0.vernier_delay_line_0.stop_strong.t67 641.061
R6805 tdc_0.vernier_delay_line_0.stop_strong.n0 tdc_0.vernier_delay_line_0.stop_strong.t78 641.061
R6806 tdc_0.vernier_delay_line_0.stop_strong.n48 tdc_0.vernier_delay_line_0.stop_strong.t41 547.874
R6807 tdc_0.vernier_delay_line_0.stop_strong.n49 tdc_0.vernier_delay_line_0.stop_strong.t54 547.874
R6808 tdc_0.vernier_delay_line_0.stop_strong.n50 tdc_0.vernier_delay_line_0.stop_strong.t32 547.874
R6809 tdc_0.vernier_delay_line_0.stop_strong.n51 tdc_0.vernier_delay_line_0.stop_strong.t34 547.874
R6810 tdc_0.vernier_delay_line_0.stop_strong.n41 tdc_0.vernier_delay_line_0.stop_strong.t65 547.874
R6811 tdc_0.vernier_delay_line_0.stop_strong.n42 tdc_0.vernier_delay_line_0.stop_strong.t85 547.874
R6812 tdc_0.vernier_delay_line_0.stop_strong.n43 tdc_0.vernier_delay_line_0.stop_strong.t50 547.874
R6813 tdc_0.vernier_delay_line_0.stop_strong.n44 tdc_0.vernier_delay_line_0.stop_strong.t63 547.874
R6814 tdc_0.vernier_delay_line_0.stop_strong.n34 tdc_0.vernier_delay_line_0.stop_strong.t83 547.874
R6815 tdc_0.vernier_delay_line_0.stop_strong.n35 tdc_0.vernier_delay_line_0.stop_strong.t47 547.874
R6816 tdc_0.vernier_delay_line_0.stop_strong.n36 tdc_0.vernier_delay_line_0.stop_strong.t62 547.874
R6817 tdc_0.vernier_delay_line_0.stop_strong.n37 tdc_0.vernier_delay_line_0.stop_strong.t84 547.874
R6818 tdc_0.vernier_delay_line_0.stop_strong.n27 tdc_0.vernier_delay_line_0.stop_strong.t42 547.874
R6819 tdc_0.vernier_delay_line_0.stop_strong.n28 tdc_0.vernier_delay_line_0.stop_strong.t44 547.874
R6820 tdc_0.vernier_delay_line_0.stop_strong.n29 tdc_0.vernier_delay_line_0.stop_strong.t57 547.874
R6821 tdc_0.vernier_delay_line_0.stop_strong.n30 tdc_0.vernier_delay_line_0.stop_strong.t73 547.874
R6822 tdc_0.vernier_delay_line_0.stop_strong.n20 tdc_0.vernier_delay_line_0.stop_strong.t53 547.874
R6823 tdc_0.vernier_delay_line_0.stop_strong.n21 tdc_0.vernier_delay_line_0.stop_strong.t69 547.874
R6824 tdc_0.vernier_delay_line_0.stop_strong.n22 tdc_0.vernier_delay_line_0.stop_strong.t71 547.874
R6825 tdc_0.vernier_delay_line_0.stop_strong.n23 tdc_0.vernier_delay_line_0.stop_strong.t36 547.874
R6826 tdc_0.vernier_delay_line_0.stop_strong.n13 tdc_0.vernier_delay_line_0.stop_strong.t68 547.874
R6827 tdc_0.vernier_delay_line_0.stop_strong.n14 tdc_0.vernier_delay_line_0.stop_strong.t35 547.874
R6828 tdc_0.vernier_delay_line_0.stop_strong.n15 tdc_0.vernier_delay_line_0.stop_strong.t51 547.874
R6829 tdc_0.vernier_delay_line_0.stop_strong.n16 tdc_0.vernier_delay_line_0.stop_strong.t64 547.874
R6830 tdc_0.vernier_delay_line_0.stop_strong.n6 tdc_0.vernier_delay_line_0.stop_strong.t33 547.874
R6831 tdc_0.vernier_delay_line_0.stop_strong.n7 tdc_0.vernier_delay_line_0.stop_strong.t60 547.874
R6832 tdc_0.vernier_delay_line_0.stop_strong.n8 tdc_0.vernier_delay_line_0.stop_strong.t82 547.874
R6833 tdc_0.vernier_delay_line_0.stop_strong.n9 tdc_0.vernier_delay_line_0.stop_strong.t46 547.874
R6834 tdc_0.vernier_delay_line_0.stop_strong.n0 tdc_0.vernier_delay_line_0.stop_strong.t43 547.874
R6835 tdc_0.vernier_delay_line_0.stop_strong.n1 tdc_0.vernier_delay_line_0.stop_strong.t55 547.874
R6836 tdc_0.vernier_delay_line_0.stop_strong.n2 tdc_0.vernier_delay_line_0.stop_strong.t72 547.874
R6837 tdc_0.vernier_delay_line_0.stop_strong.n3 tdc_0.vernier_delay_line_0.stop_strong.t37 547.874
R6838 tdc_0.vernier_delay_line_0.stop_strong.n53 tdc_0.vernier_delay_line_0.stop_strong.n51 189.41
R6839 tdc_0.vernier_delay_line_0.stop_strong.n46 tdc_0.vernier_delay_line_0.stop_strong.n44 189.41
R6840 tdc_0.vernier_delay_line_0.stop_strong.n39 tdc_0.vernier_delay_line_0.stop_strong.n37 189.41
R6841 tdc_0.vernier_delay_line_0.stop_strong.n32 tdc_0.vernier_delay_line_0.stop_strong.n30 189.41
R6842 tdc_0.vernier_delay_line_0.stop_strong.n25 tdc_0.vernier_delay_line_0.stop_strong.n23 189.41
R6843 tdc_0.vernier_delay_line_0.stop_strong.n18 tdc_0.vernier_delay_line_0.stop_strong.n16 189.41
R6844 tdc_0.vernier_delay_line_0.stop_strong.n11 tdc_0.vernier_delay_line_0.stop_strong.n9 189.41
R6845 tdc_0.vernier_delay_line_0.stop_strong.n5 tdc_0.vernier_delay_line_0.stop_strong.n3 189.41
R6846 tdc_0.vernier_delay_line_0.stop_strong.n49 tdc_0.vernier_delay_line_0.stop_strong.n48 93.1872
R6847 tdc_0.vernier_delay_line_0.stop_strong.n50 tdc_0.vernier_delay_line_0.stop_strong.n49 93.1872
R6848 tdc_0.vernier_delay_line_0.stop_strong.n51 tdc_0.vernier_delay_line_0.stop_strong.n50 93.1872
R6849 tdc_0.vernier_delay_line_0.stop_strong.n42 tdc_0.vernier_delay_line_0.stop_strong.n41 93.1872
R6850 tdc_0.vernier_delay_line_0.stop_strong.n43 tdc_0.vernier_delay_line_0.stop_strong.n42 93.1872
R6851 tdc_0.vernier_delay_line_0.stop_strong.n44 tdc_0.vernier_delay_line_0.stop_strong.n43 93.1872
R6852 tdc_0.vernier_delay_line_0.stop_strong.n35 tdc_0.vernier_delay_line_0.stop_strong.n34 93.1872
R6853 tdc_0.vernier_delay_line_0.stop_strong.n36 tdc_0.vernier_delay_line_0.stop_strong.n35 93.1872
R6854 tdc_0.vernier_delay_line_0.stop_strong.n37 tdc_0.vernier_delay_line_0.stop_strong.n36 93.1872
R6855 tdc_0.vernier_delay_line_0.stop_strong.n28 tdc_0.vernier_delay_line_0.stop_strong.n27 93.1872
R6856 tdc_0.vernier_delay_line_0.stop_strong.n29 tdc_0.vernier_delay_line_0.stop_strong.n28 93.1872
R6857 tdc_0.vernier_delay_line_0.stop_strong.n30 tdc_0.vernier_delay_line_0.stop_strong.n29 93.1872
R6858 tdc_0.vernier_delay_line_0.stop_strong.n21 tdc_0.vernier_delay_line_0.stop_strong.n20 93.1872
R6859 tdc_0.vernier_delay_line_0.stop_strong.n22 tdc_0.vernier_delay_line_0.stop_strong.n21 93.1872
R6860 tdc_0.vernier_delay_line_0.stop_strong.n23 tdc_0.vernier_delay_line_0.stop_strong.n22 93.1872
R6861 tdc_0.vernier_delay_line_0.stop_strong.n14 tdc_0.vernier_delay_line_0.stop_strong.n13 93.1872
R6862 tdc_0.vernier_delay_line_0.stop_strong.n15 tdc_0.vernier_delay_line_0.stop_strong.n14 93.1872
R6863 tdc_0.vernier_delay_line_0.stop_strong.n16 tdc_0.vernier_delay_line_0.stop_strong.n15 93.1872
R6864 tdc_0.vernier_delay_line_0.stop_strong.n7 tdc_0.vernier_delay_line_0.stop_strong.n6 93.1872
R6865 tdc_0.vernier_delay_line_0.stop_strong.n8 tdc_0.vernier_delay_line_0.stop_strong.n7 93.1872
R6866 tdc_0.vernier_delay_line_0.stop_strong.n9 tdc_0.vernier_delay_line_0.stop_strong.n8 93.1872
R6867 tdc_0.vernier_delay_line_0.stop_strong.n1 tdc_0.vernier_delay_line_0.stop_strong.n0 93.1872
R6868 tdc_0.vernier_delay_line_0.stop_strong.n2 tdc_0.vernier_delay_line_0.stop_strong.n1 93.1872
R6869 tdc_0.vernier_delay_line_0.stop_strong.n3 tdc_0.vernier_delay_line_0.stop_strong.n2 93.1872
R6870 tdc_0.vernier_delay_line_0.stop_strong.n82 tdc_0.vernier_delay_line_0.stop_strong.t21 85.2499
R6871 tdc_0.vernier_delay_line_0.stop_strong.n80 tdc_0.vernier_delay_line_0.stop_strong.t28 85.2499
R6872 tdc_0.vernier_delay_line_0.stop_strong.n78 tdc_0.vernier_delay_line_0.stop_strong.t18 85.2499
R6873 tdc_0.vernier_delay_line_0.stop_strong.n76 tdc_0.vernier_delay_line_0.stop_strong.t24 85.2499
R6874 tdc_0.vernier_delay_line_0.stop_strong.n74 tdc_0.vernier_delay_line_0.stop_strong.t22 85.2499
R6875 tdc_0.vernier_delay_line_0.stop_strong.n72 tdc_0.vernier_delay_line_0.stop_strong.t29 85.2499
R6876 tdc_0.vernier_delay_line_0.stop_strong.n70 tdc_0.vernier_delay_line_0.stop_strong.t19 85.2499
R6877 tdc_0.vernier_delay_line_0.stop_strong.n68 tdc_0.vernier_delay_line_0.stop_strong.t25 85.2499
R6878 tdc_0.vernier_delay_line_0.stop_strong.n66 tdc_0.vernier_delay_line_0.stop_strong.t16 85.2499
R6879 tdc_0.vernier_delay_line_0.stop_strong.n64 tdc_0.vernier_delay_line_0.stop_strong.t26 85.2499
R6880 tdc_0.vernier_delay_line_0.stop_strong.n62 tdc_0.vernier_delay_line_0.stop_strong.t17 85.2499
R6881 tdc_0.vernier_delay_line_0.stop_strong.n60 tdc_0.vernier_delay_line_0.stop_strong.t23 85.2499
R6882 tdc_0.vernier_delay_line_0.stop_strong.n58 tdc_0.vernier_delay_line_0.stop_strong.t30 85.2499
R6883 tdc_0.vernier_delay_line_0.stop_strong.n56 tdc_0.vernier_delay_line_0.stop_strong.t20 85.2499
R6884 tdc_0.vernier_delay_line_0.stop_strong.n55 tdc_0.vernier_delay_line_0.stop_strong.t27 85.2499
R6885 tdc_0.vernier_delay_line_0.stop_strong.n86 tdc_0.vernier_delay_line_0.stop_strong.t31 84.7281
R6886 tdc_0.vernier_delay_line_0.stop_strong.n85 tdc_0.vernier_delay_line_0.stop_strong.t1 83.7172
R6887 tdc_0.vernier_delay_line_0.stop_strong.n82 tdc_0.vernier_delay_line_0.stop_strong.t7 83.7172
R6888 tdc_0.vernier_delay_line_0.stop_strong.n80 tdc_0.vernier_delay_line_0.stop_strong.t14 83.7172
R6889 tdc_0.vernier_delay_line_0.stop_strong.n78 tdc_0.vernier_delay_line_0.stop_strong.t4 83.7172
R6890 tdc_0.vernier_delay_line_0.stop_strong.n76 tdc_0.vernier_delay_line_0.stop_strong.t10 83.7172
R6891 tdc_0.vernier_delay_line_0.stop_strong.n74 tdc_0.vernier_delay_line_0.stop_strong.t8 83.7172
R6892 tdc_0.vernier_delay_line_0.stop_strong.n72 tdc_0.vernier_delay_line_0.stop_strong.t15 83.7172
R6893 tdc_0.vernier_delay_line_0.stop_strong.n70 tdc_0.vernier_delay_line_0.stop_strong.t5 83.7172
R6894 tdc_0.vernier_delay_line_0.stop_strong.n68 tdc_0.vernier_delay_line_0.stop_strong.t11 83.7172
R6895 tdc_0.vernier_delay_line_0.stop_strong.n66 tdc_0.vernier_delay_line_0.stop_strong.t2 83.7172
R6896 tdc_0.vernier_delay_line_0.stop_strong.n64 tdc_0.vernier_delay_line_0.stop_strong.t12 83.7172
R6897 tdc_0.vernier_delay_line_0.stop_strong.n62 tdc_0.vernier_delay_line_0.stop_strong.t3 83.7172
R6898 tdc_0.vernier_delay_line_0.stop_strong.n60 tdc_0.vernier_delay_line_0.stop_strong.t9 83.7172
R6899 tdc_0.vernier_delay_line_0.stop_strong.n58 tdc_0.vernier_delay_line_0.stop_strong.t0 83.7172
R6900 tdc_0.vernier_delay_line_0.stop_strong.n56 tdc_0.vernier_delay_line_0.stop_strong.t6 83.7172
R6901 tdc_0.vernier_delay_line_0.stop_strong.n55 tdc_0.vernier_delay_line_0.stop_strong.t13 83.7172
R6902 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n5 11.8482
R6903 tdc_0.vernier_delay_line_0.stop_strong.n54 tdc_0.vernier_delay_line_0.stop_strong.n53 9.66066
R6904 tdc_0.vernier_delay_line_0.stop_strong.n47 tdc_0.vernier_delay_line_0.stop_strong.n46 9.66066
R6905 tdc_0.vernier_delay_line_0.stop_strong.n40 tdc_0.vernier_delay_line_0.stop_strong.n39 9.66066
R6906 tdc_0.vernier_delay_line_0.stop_strong.n33 tdc_0.vernier_delay_line_0.stop_strong.n32 9.66066
R6907 tdc_0.vernier_delay_line_0.stop_strong.n26 tdc_0.vernier_delay_line_0.stop_strong.n25 9.66066
R6908 tdc_0.vernier_delay_line_0.stop_strong.n19 tdc_0.vernier_delay_line_0.stop_strong.n18 9.66066
R6909 tdc_0.vernier_delay_line_0.stop_strong.n12 tdc_0.vernier_delay_line_0.stop_strong.n11 9.66066
R6910 tdc_0.vernier_delay_line_0.stop_strong.n84 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk 8.04701
R6911 tdc_0.vernier_delay_line_0.stop_strong.n57 tdc_0.vernier_delay_line_0.stop_strong.n55 5.16238
R6912 tdc_0.vernier_delay_line_0.stop_strong.n83 tdc_0.vernier_delay_line_0.stop_strong.n82 4.64452
R6913 tdc_0.vernier_delay_line_0.stop_strong.n81 tdc_0.vernier_delay_line_0.stop_strong.n80 4.64452
R6914 tdc_0.vernier_delay_line_0.stop_strong.n79 tdc_0.vernier_delay_line_0.stop_strong.n78 4.64452
R6915 tdc_0.vernier_delay_line_0.stop_strong.n77 tdc_0.vernier_delay_line_0.stop_strong.n76 4.64452
R6916 tdc_0.vernier_delay_line_0.stop_strong.n75 tdc_0.vernier_delay_line_0.stop_strong.n74 4.64452
R6917 tdc_0.vernier_delay_line_0.stop_strong.n73 tdc_0.vernier_delay_line_0.stop_strong.n72 4.64452
R6918 tdc_0.vernier_delay_line_0.stop_strong.n71 tdc_0.vernier_delay_line_0.stop_strong.n70 4.64452
R6919 tdc_0.vernier_delay_line_0.stop_strong.n69 tdc_0.vernier_delay_line_0.stop_strong.n68 4.64452
R6920 tdc_0.vernier_delay_line_0.stop_strong.n67 tdc_0.vernier_delay_line_0.stop_strong.n66 4.64452
R6921 tdc_0.vernier_delay_line_0.stop_strong.n65 tdc_0.vernier_delay_line_0.stop_strong.n64 4.64452
R6922 tdc_0.vernier_delay_line_0.stop_strong.n63 tdc_0.vernier_delay_line_0.stop_strong.n62 4.64452
R6923 tdc_0.vernier_delay_line_0.stop_strong.n61 tdc_0.vernier_delay_line_0.stop_strong.n60 4.64452
R6924 tdc_0.vernier_delay_line_0.stop_strong.n59 tdc_0.vernier_delay_line_0.stop_strong.n58 4.64452
R6925 tdc_0.vernier_delay_line_0.stop_strong.n57 tdc_0.vernier_delay_line_0.stop_strong.n56 4.64452
R6926 tdc_0.vernier_delay_line_0.stop_strong.n85 tdc_0.vernier_delay_line_0.stop_strong.n84 4.64452
R6927 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n12 2.188
R6928 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n19 2.188
R6929 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n26 2.188
R6930 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n33 2.188
R6931 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n40 2.188
R6932 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n47 2.188
R6933 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n54 2.188
R6934 tdc_0.vernier_delay_line_0.stop_strong.n53 tdc_0.vernier_delay_line_0.stop_strong.n52 1.05649
R6935 tdc_0.vernier_delay_line_0.stop_strong.n46 tdc_0.vernier_delay_line_0.stop_strong.n45 1.05649
R6936 tdc_0.vernier_delay_line_0.stop_strong.n39 tdc_0.vernier_delay_line_0.stop_strong.n38 1.05649
R6937 tdc_0.vernier_delay_line_0.stop_strong.n32 tdc_0.vernier_delay_line_0.stop_strong.n31 1.05649
R6938 tdc_0.vernier_delay_line_0.stop_strong.n25 tdc_0.vernier_delay_line_0.stop_strong.n24 1.05649
R6939 tdc_0.vernier_delay_line_0.stop_strong.n18 tdc_0.vernier_delay_line_0.stop_strong.n17 1.05649
R6940 tdc_0.vernier_delay_line_0.stop_strong.n11 tdc_0.vernier_delay_line_0.stop_strong.n10 1.05649
R6941 tdc_0.vernier_delay_line_0.stop_strong.n5 tdc_0.vernier_delay_line_0.stop_strong.n4 1.05649
R6942 tdc_0.vernier_delay_line_0.stop_strong.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk 0.6655
R6943 tdc_0.vernier_delay_line_0.stop_strong.n19 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk 0.6655
R6944 tdc_0.vernier_delay_line_0.stop_strong.n26 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk 0.6655
R6945 tdc_0.vernier_delay_line_0.stop_strong.n33 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk 0.6655
R6946 tdc_0.vernier_delay_line_0.stop_strong.n40 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk 0.6655
R6947 tdc_0.vernier_delay_line_0.stop_strong.n47 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk 0.6655
R6948 tdc_0.vernier_delay_line_0.stop_strong.n54 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk 0.6655
R6949 tdc_0.vernier_delay_line_0.stop_strong.n83 tdc_0.vernier_delay_line_0.stop_strong.n81 0.518357
R6950 tdc_0.vernier_delay_line_0.stop_strong.n81 tdc_0.vernier_delay_line_0.stop_strong.n79 0.518357
R6951 tdc_0.vernier_delay_line_0.stop_strong.n79 tdc_0.vernier_delay_line_0.stop_strong.n77 0.518357
R6952 tdc_0.vernier_delay_line_0.stop_strong.n77 tdc_0.vernier_delay_line_0.stop_strong.n75 0.518357
R6953 tdc_0.vernier_delay_line_0.stop_strong.n75 tdc_0.vernier_delay_line_0.stop_strong.n73 0.518357
R6954 tdc_0.vernier_delay_line_0.stop_strong.n73 tdc_0.vernier_delay_line_0.stop_strong.n71 0.518357
R6955 tdc_0.vernier_delay_line_0.stop_strong.n71 tdc_0.vernier_delay_line_0.stop_strong.n69 0.518357
R6956 tdc_0.vernier_delay_line_0.stop_strong.n69 tdc_0.vernier_delay_line_0.stop_strong.n67 0.518357
R6957 tdc_0.vernier_delay_line_0.stop_strong.n67 tdc_0.vernier_delay_line_0.stop_strong.n65 0.518357
R6958 tdc_0.vernier_delay_line_0.stop_strong.n65 tdc_0.vernier_delay_line_0.stop_strong.n63 0.518357
R6959 tdc_0.vernier_delay_line_0.stop_strong.n63 tdc_0.vernier_delay_line_0.stop_strong.n61 0.518357
R6960 tdc_0.vernier_delay_line_0.stop_strong.n61 tdc_0.vernier_delay_line_0.stop_strong.n59 0.518357
R6961 tdc_0.vernier_delay_line_0.stop_strong.n59 tdc_0.vernier_delay_line_0.stop_strong.n57 0.518357
R6962 tdc_0.vernier_delay_line_0.stop_strong.n84 tdc_0.vernier_delay_line_0.stop_strong.n83 0.497131
R6963 tdc_0.vernier_delay_line_0.stop_strong.n86 tdc_0.vernier_delay_line_0.stop_strong.n85 0.3755
R6964 tdc_0.stop_buffer_0.stop_strong tdc_0.vernier_delay_line_0.stop_strong.n86 0.234296
R6965 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 784.053
R6966 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 784.053
R6967 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 784.053
R6968 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 784.053
R6969 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 539.841
R6970 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 539.841
R6971 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 539.841
R6972 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 539.841
R6973 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 215.293
R6974 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 215.293
R6975 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 215.293
R6976 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 215.293
R6977 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 168.659
R6978 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 167.992
R6979 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 166.144
R6980 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 165.8
R6981 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 85.2499
R6982 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 85.2499
R6983 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 83.7172
R6984 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 83.7172
R6985 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 75.7282
R6986 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 66.3172
R6987 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 36.1505
R6988 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 36.1505
R6989 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 34.5438
R6990 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 34.5438
R6991 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 17.4005
R6992 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 17.4005
R6993 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 17.2391
R6994 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 9.52217
R6995 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 9.52217
R6996 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 6.39571
R6997 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 5.30824
R6998 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 4.94887
R6999 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 1.64112
R7000 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 1.06691
R7001 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd 0.930188
R7002 a_10108_39954.n2 a_10108_39954.n1 34.9195
R7003 a_10108_39954.n3 a_10108_39954.n2 25.5407
R7004 a_10108_39954.n2 a_10108_39954.n0 25.2907
R7005 a_10108_39954.n1 a_10108_39954.t4 5.8005
R7006 a_10108_39954.n1 a_10108_39954.t5 5.8005
R7007 a_10108_39954.n0 a_10108_39954.t3 5.8005
R7008 a_10108_39954.n0 a_10108_39954.t2 5.8005
R7009 a_10108_39954.t0 a_10108_39954.n3 5.8005
R7010 a_10108_39954.n3 a_10108_39954.t1 5.8005
R7011 a_10958_39338.n1 a_10958_39338.t0 31.9657
R7012 a_10958_39338.n1 a_10958_39338.n0 25.8125
R7013 a_10958_39338.n3 a_10958_39338.n2 25.8125
R7014 a_10958_39338.n5 a_10958_39338.n4 25.8125
R7015 a_10958_39338.n10 a_10958_39338.n9 25.7038
R7016 a_10958_39338.n9 a_10958_39338.n8 25.3505
R7017 a_10958_39338.n7 a_10958_39338.n6 24.288
R7018 a_10958_39338.n6 a_10958_39338.t3 5.8005
R7019 a_10958_39338.n6 a_10958_39338.t10 5.8005
R7020 a_10958_39338.n0 a_10958_39338.t8 5.8005
R7021 a_10958_39338.n0 a_10958_39338.t2 5.8005
R7022 a_10958_39338.n2 a_10958_39338.t1 5.8005
R7023 a_10958_39338.n2 a_10958_39338.t11 5.8005
R7024 a_10958_39338.n4 a_10958_39338.t9 5.8005
R7025 a_10958_39338.n4 a_10958_39338.t12 5.8005
R7026 a_10958_39338.n8 a_10958_39338.t5 5.8005
R7027 a_10958_39338.n8 a_10958_39338.t6 5.8005
R7028 a_10958_39338.t7 a_10958_39338.n10 5.8005
R7029 a_10958_39338.n10 a_10958_39338.t4 5.8005
R7030 a_10958_39338.n7 a_10958_39338.n5 1.87822
R7031 a_10958_39338.n9 a_10958_39338.n7 1.41626
R7032 a_10958_39338.n3 a_10958_39338.n1 0.353761
R7033 a_10958_39338.n5 a_10958_39338.n3 0.353761
R7034 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 890.727
R7035 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 742.783
R7036 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 641.061
R7037 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7038 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7039 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7040 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7041 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7042 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7043 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7044 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7045 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R7046 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R7047 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R7048 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7049 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 8.91506
R7050 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7051 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7052 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7053 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7054 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 879.481
R7055 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 742.783
R7056 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 641.061
R7057 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 623.388
R7058 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 547.874
R7059 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 431.807
R7060 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 427.875
R7061 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 333.161
R7062 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7063 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 168.077
R7064 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R7065 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7066 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7067 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 11.1806
R7068 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7069 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7070 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R7071 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7072 a_10108_28544.n2 a_10108_28544.n1 34.9195
R7073 a_10108_28544.n3 a_10108_28544.n2 25.5407
R7074 a_10108_28544.n2 a_10108_28544.n0 25.2907
R7075 a_10108_28544.n1 a_10108_28544.t3 5.8005
R7076 a_10108_28544.n1 a_10108_28544.t4 5.8005
R7077 a_10108_28544.n0 a_10108_28544.t5 5.8005
R7078 a_10108_28544.n0 a_10108_28544.t2 5.8005
R7079 a_10108_28544.n3 a_10108_28544.t0 5.8005
R7080 a_10108_28544.t1 a_10108_28544.n3 5.8005
R7081 a_10958_23364.n1 a_10958_23364.t1 31.9657
R7082 a_10958_23364.n1 a_10958_23364.n0 25.8125
R7083 a_10958_23364.n3 a_10958_23364.n2 25.8125
R7084 a_10958_23364.n5 a_10958_23364.n4 25.8125
R7085 a_10958_23364.n10 a_10958_23364.n9 25.7038
R7086 a_10958_23364.n9 a_10958_23364.n8 25.3505
R7087 a_10958_23364.n7 a_10958_23364.n6 24.288
R7088 a_10958_23364.n6 a_10958_23364.t3 5.8005
R7089 a_10958_23364.n6 a_10958_23364.t11 5.8005
R7090 a_10958_23364.n0 a_10958_23364.t9 5.8005
R7091 a_10958_23364.n0 a_10958_23364.t2 5.8005
R7092 a_10958_23364.n2 a_10958_23364.t0 5.8005
R7093 a_10958_23364.n2 a_10958_23364.t10 5.8005
R7094 a_10958_23364.n4 a_10958_23364.t12 5.8005
R7095 a_10958_23364.n4 a_10958_23364.t8 5.8005
R7096 a_10958_23364.n8 a_10958_23364.t4 5.8005
R7097 a_10958_23364.n8 a_10958_23364.t5 5.8005
R7098 a_10958_23364.n10 a_10958_23364.t6 5.8005
R7099 a_10958_23364.t7 a_10958_23364.n10 5.8005
R7100 a_10958_23364.n7 a_10958_23364.n5 1.87822
R7101 a_10958_23364.n9 a_10958_23364.n7 1.41626
R7102 a_10958_23364.n3 a_10958_23364.n1 0.353761
R7103 a_10958_23364.n5 a_10958_23364.n3 0.353761
R7104 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 628.097
R7105 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 622.766
R7106 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 523.774
R7107 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 304.647
R7108 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 304.647
R7109 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 202.44
R7110 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 169.062
R7111 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 166.237
R7112 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R7113 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R7114 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R7115 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 5.48979
R7116 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 4.5005
R7117 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 1.09595
R7118 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 879.481
R7119 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7120 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 641.061
R7121 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 623.388
R7122 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 547.874
R7123 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 431.807
R7124 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 427.875
R7125 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7126 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7127 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7128 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7129 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 31.2972
R7130 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7131 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 11.1806
R7132 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7133 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R7134 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R7135 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7136 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 890.727
R7137 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 742.783
R7138 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 641.061
R7139 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 623.388
R7140 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7141 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7142 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7143 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7144 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7145 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7146 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7147 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R7148 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R7149 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R7150 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7151 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 8.91506
R7152 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7153 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7154 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7155 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7156 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 879.481
R7157 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 742.783
R7158 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 641.061
R7159 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 623.388
R7160 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 547.874
R7161 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 431.807
R7162 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 427.875
R7163 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7164 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7165 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7166 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7167 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R7168 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7169 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 11.1806
R7170 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7171 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R7172 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7173 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7174 a_10108_35390.n2 a_10108_35390.n1 34.9195
R7175 a_10108_35390.n3 a_10108_35390.n2 25.5407
R7176 a_10108_35390.n2 a_10108_35390.n0 25.2907
R7177 a_10108_35390.n1 a_10108_35390.t4 5.8005
R7178 a_10108_35390.n1 a_10108_35390.t5 5.8005
R7179 a_10108_35390.n0 a_10108_35390.t3 5.8005
R7180 a_10108_35390.n0 a_10108_35390.t0 5.8005
R7181 a_10108_35390.n3 a_10108_35390.t1 5.8005
R7182 a_10108_35390.t2 a_10108_35390.n3 5.8005
R7183 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 879.481
R7184 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7185 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 641.061
R7186 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 623.388
R7187 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 547.874
R7188 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 431.807
R7189 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 427.875
R7190 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7191 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7192 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7193 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7194 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R7195 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7196 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 11.1806
R7197 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7198 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7199 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R7200 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7201 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 890.727
R7202 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 742.783
R7203 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 641.061
R7204 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7205 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7206 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 431.807
R7207 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7208 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7209 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7210 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7211 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7212 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R7213 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R7214 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R7215 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7216 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 8.91506
R7217 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7218 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7219 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7220 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7221 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 628.097
R7222 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 622.766
R7223 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 523.774
R7224 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 304.647
R7225 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 304.647
R7226 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 202.44
R7227 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 169.062
R7228 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 166.237
R7229 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 84.7557
R7230 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 84.1197
R7231 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 12.6535
R7232 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 5.48979
R7233 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 4.5005
R7234 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 1.09595
R7235 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 552.84
R7236 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 552.84
R7237 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 552.84
R7238 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 552.84
R7239 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 539.841
R7240 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 539.841
R7241 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 539.841
R7242 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 539.841
R7243 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 215.293
R7244 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 215.293
R7245 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 215.293
R7246 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 215.293
R7247 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 166.468
R7248 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 166.149
R7249 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 165.8
R7250 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 165.8
R7251 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 85.1574
R7252 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 83.8097
R7253 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 83.8097
R7254 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 83.7172
R7255 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 74.288
R7256 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 67.7574
R7257 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 36.1505
R7258 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 36.1505
R7259 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 34.5438
R7260 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 34.5438
R7261 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 17.4005
R7262 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 17.4005
R7263 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 16.09
R7264 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 11.8364
R7265 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 9.52217
R7266 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 9.52217
R7267 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d 5.96628
R7268 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 5.83219
R7269 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 5.74235
R7270 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 5.49235
R7271 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 2.48878
R7272 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 1.44072
R7273 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 1.32081
R7274 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 628.097
R7275 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 622.766
R7276 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 523.774
R7277 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 304.647
R7278 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 304.647
R7279 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 202.44
R7280 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 169.062
R7281 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 166.237
R7282 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 84.7557
R7283 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 84.1197
R7284 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 12.6535
R7285 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 5.48979
R7286 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 4.5005
R7287 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 1.09595
R7288 a_10958_37056.n2 a_10958_37056.t11 31.9657
R7289 a_10958_37056.n2 a_10958_37056.n1 25.8125
R7290 a_10958_37056.n4 a_10958_37056.n3 25.8125
R7291 a_10958_37056.n6 a_10958_37056.n5 25.8125
R7292 a_10958_37056.n9 a_10958_37056.n0 25.7038
R7293 a_10958_37056.n10 a_10958_37056.n9 25.3505
R7294 a_10958_37056.n8 a_10958_37056.n7 24.288
R7295 a_10958_37056.n7 a_10958_37056.t5 5.8005
R7296 a_10958_37056.n7 a_10958_37056.t3 5.8005
R7297 a_10958_37056.n1 a_10958_37056.t0 5.8005
R7298 a_10958_37056.n1 a_10958_37056.t10 5.8005
R7299 a_10958_37056.n3 a_10958_37056.t12 5.8005
R7300 a_10958_37056.n3 a_10958_37056.t1 5.8005
R7301 a_10958_37056.n5 a_10958_37056.t9 5.8005
R7302 a_10958_37056.n5 a_10958_37056.t2 5.8005
R7303 a_10958_37056.n0 a_10958_37056.t7 5.8005
R7304 a_10958_37056.n0 a_10958_37056.t4 5.8005
R7305 a_10958_37056.n10 a_10958_37056.t6 5.8005
R7306 a_10958_37056.t8 a_10958_37056.n10 5.8005
R7307 a_10958_37056.n8 a_10958_37056.n6 1.87822
R7308 a_10958_37056.n9 a_10958_37056.n8 1.41626
R7309 a_10958_37056.n4 a_10958_37056.n2 0.353761
R7310 a_10958_37056.n6 a_10958_37056.n4 0.353761
R7311 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 890.727
R7312 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 742.783
R7313 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 641.061
R7314 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 623.388
R7315 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 547.874
R7316 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 431.807
R7317 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 427.875
R7318 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7319 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7320 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7321 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7322 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 31.2103
R7323 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R7324 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R7325 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7326 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 8.91506
R7327 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7328 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7329 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7330 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7331 a_10108_26262.n2 a_10108_26262.n1 34.9195
R7332 a_10108_26262.n3 a_10108_26262.n2 25.5407
R7333 a_10108_26262.n2 a_10108_26262.n0 25.2907
R7334 a_10108_26262.n1 a_10108_26262.t4 5.8005
R7335 a_10108_26262.n1 a_10108_26262.t0 5.8005
R7336 a_10108_26262.n0 a_10108_26262.t3 5.8005
R7337 a_10108_26262.n0 a_10108_26262.t5 5.8005
R7338 a_10108_26262.t2 a_10108_26262.n3 5.8005
R7339 a_10108_26262.n3 a_10108_26262.t1 5.8005
R7340 uo_out[6].n0 uo_out[6].t5 734.539
R7341 uo_out[6].n0 uo_out[6].t4 233.26
R7342 uo_out[6].n2 uo_out[6].n0 162.335
R7343 uo_out[6].n2 uo_out[6].n1 75.5733
R7344 uo_out[6].n4 uo_out[6].n3 66.3172
R7345 uo_out[6].n3 uo_out[6].t3 17.4005
R7346 uo_out[6].n3 uo_out[6].t0 17.4005
R7347 uo_out[6].n5 uo_out[6] 16.4025
R7348 uo_out[6].n1 uo_out[6].t1 9.52217
R7349 uo_out[6].n1 uo_out[6].t2 9.52217
R7350 uo_out[6].n5 uo_out[6].n4 5.02496
R7351 uo_out[6].n4 uo_out[6].n2 0.438
R7352 uo_out[6] uo_out[6].n5 0.063
R7353 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 628.097
R7354 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 622.766
R7355 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 523.774
R7356 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 304.647
R7357 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 304.647
R7358 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 202.44
R7359 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 169.062
R7360 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 166.237
R7361 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 84.7557
R7362 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 84.1197
R7363 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 12.6535
R7364 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 5.48979
R7365 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 4.5005
R7366 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 1.09595
R7367 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 539.841
R7368 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 539.841
R7369 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 539.841
R7370 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 539.841
R7371 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 215.293
R7372 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 215.293
R7373 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 215.293
R7374 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 215.293
R7375 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 166.144
R7376 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 165.8
R7377 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 85.2499
R7378 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 85.2499
R7379 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 83.7172
R7380 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 83.7172
R7381 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 75.7282
R7382 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 66.3172
R7383 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 36.1505
R7384 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 36.1505
R7385 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 34.5438
R7386 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 34.5438
R7387 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 17.4005
R7388 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 17.4005
R7389 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 9.52217
R7390 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 9.52217
R7391 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 6.39571
R7392 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 5.30824
R7393 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 4.94887
R7394 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 1.06691
R7395 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 0.160656
R7396 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 539.841
R7397 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 539.841
R7398 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 539.841
R7399 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 539.841
R7400 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 215.293
R7401 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 215.293
R7402 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 215.293
R7403 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 215.293
R7404 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 166.149
R7405 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 165.8
R7406 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 85.1574
R7407 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 85.1574
R7408 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 83.8097
R7409 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 83.8097
R7410 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 74.288
R7411 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 67.7574
R7412 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 36.1505
R7413 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 36.1505
R7414 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 34.5438
R7415 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 34.5438
R7416 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 17.4005
R7417 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 17.4005
R7418 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 11.8364
R7419 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 9.52217
R7420 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 9.52217
R7421 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 5.83219
R7422 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 5.74235
R7423 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 5.49235
R7424 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 1.32081
R7425 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 0.285656
R7426 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 539.841
R7427 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 539.841
R7428 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 539.841
R7429 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 539.841
R7430 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 215.293
R7431 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 215.293
R7432 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 215.293
R7433 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 215.293
R7434 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 166.144
R7435 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 165.8
R7436 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 85.2499
R7437 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 85.2499
R7438 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 83.7172
R7439 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 83.7172
R7440 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 75.7282
R7441 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 66.3172
R7442 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 36.1505
R7443 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 36.1505
R7444 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 34.5438
R7445 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 34.5438
R7446 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 17.4005
R7447 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 17.4005
R7448 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 9.52217
R7449 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 9.52217
R7450 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 6.39571
R7451 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 5.30824
R7452 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 4.94887
R7453 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 1.41456
R7454 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 539.841
R7455 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 539.841
R7456 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 539.841
R7457 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 539.841
R7458 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 215.293
R7459 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 215.293
R7460 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 215.293
R7461 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 215.293
R7462 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 166.149
R7463 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 165.8
R7464 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 85.1574
R7465 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 85.1574
R7466 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 83.8097
R7467 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 83.8097
R7468 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 74.288
R7469 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 67.7574
R7470 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 36.1505
R7471 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 36.1505
R7472 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 34.5438
R7473 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 34.5438
R7474 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 17.4005
R7475 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 17.4005
R7476 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 11.8364
R7477 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 9.52217
R7478 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 9.52217
R7479 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 5.83219
R7480 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 5.74235
R7481 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 5.49235
R7482 tdc_0.diff_gen_0.delay_unit_2_4.out_1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 1.32081
R7483 tdc_0.diff_gen_0.delay_unit_2_4.out_1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 0.53175
R7484 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 552.84
R7485 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 552.84
R7486 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 552.84
R7487 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 552.84
R7488 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 539.841
R7489 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 539.841
R7490 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 539.841
R7491 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 539.841
R7492 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 215.293
R7493 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 215.293
R7494 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 215.293
R7495 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 215.293
R7496 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 166.468
R7497 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 166.149
R7498 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 165.8
R7499 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 165.8
R7500 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 85.1574
R7501 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 83.8097
R7502 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 83.8097
R7503 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 83.7172
R7504 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 74.288
R7505 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 67.7574
R7506 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 36.1505
R7507 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 36.1505
R7508 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 34.5438
R7509 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 34.5438
R7510 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 17.4005
R7511 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 17.4005
R7512 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 16.09
R7513 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 11.8364
R7514 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 9.52217
R7515 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 9.52217
R7516 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 5.96628
R7517 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 5.83219
R7518 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 5.74235
R7519 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 5.49235
R7520 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 1.44072
R7521 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.32081
R7522 a_10958_34774.n2 a_10958_34774.t12 31.9657
R7523 a_10958_34774.n2 a_10958_34774.n1 25.8125
R7524 a_10958_34774.n4 a_10958_34774.n3 25.8125
R7525 a_10958_34774.n6 a_10958_34774.n5 25.8125
R7526 a_10958_34774.n9 a_10958_34774.n0 25.7038
R7527 a_10958_34774.n10 a_10958_34774.n9 25.3505
R7528 a_10958_34774.n8 a_10958_34774.n7 24.288
R7529 a_10958_34774.n7 a_10958_34774.t6 5.8005
R7530 a_10958_34774.n7 a_10958_34774.t9 5.8005
R7531 a_10958_34774.n1 a_10958_34774.t11 5.8005
R7532 a_10958_34774.n1 a_10958_34774.t2 5.8005
R7533 a_10958_34774.n3 a_10958_34774.t1 5.8005
R7534 a_10958_34774.n3 a_10958_34774.t10 5.8005
R7535 a_10958_34774.n5 a_10958_34774.t3 5.8005
R7536 a_10958_34774.n5 a_10958_34774.t0 5.8005
R7537 a_10958_34774.n0 a_10958_34774.t5 5.8005
R7538 a_10958_34774.n0 a_10958_34774.t7 5.8005
R7539 a_10958_34774.t8 a_10958_34774.n10 5.8005
R7540 a_10958_34774.n10 a_10958_34774.t4 5.8005
R7541 a_10958_34774.n8 a_10958_34774.n6 1.87822
R7542 a_10958_34774.n9 a_10958_34774.n8 1.41626
R7543 a_10958_34774.n4 a_10958_34774.n2 0.353761
R7544 a_10958_34774.n6 a_10958_34774.n4 0.353761
R7545 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 539.841
R7546 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 539.841
R7547 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 539.841
R7548 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 539.841
R7549 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 215.293
R7550 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 215.293
R7551 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 215.293
R7552 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 215.293
R7553 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 166.144
R7554 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 165.8
R7555 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 85.2499
R7556 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 85.2499
R7557 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 83.7172
R7558 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 83.7172
R7559 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 75.7282
R7560 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 66.3172
R7561 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 36.1505
R7562 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 36.1505
R7563 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 34.5438
R7564 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 34.5438
R7565 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 17.4005
R7566 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 17.4005
R7567 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 9.52217
R7568 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 9.52217
R7569 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 6.39571
R7570 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 5.30824
R7571 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 4.94887
R7572 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 1.41456
R7573 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 784.053
R7574 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 784.053
R7575 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 784.053
R7576 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 784.053
R7577 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 539.841
R7578 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 539.841
R7579 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 539.841
R7580 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 539.841
R7581 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 215.293
R7582 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 215.293
R7583 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 215.293
R7584 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 215.293
R7585 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 168.659
R7586 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 167.992
R7587 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 166.144
R7588 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 165.8
R7589 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 85.2499
R7590 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 85.2499
R7591 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 83.7172
R7592 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 83.7172
R7593 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 75.7282
R7594 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 66.3172
R7595 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 36.1505
R7596 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 36.1505
R7597 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 34.5438
R7598 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 34.5438
R7599 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 17.4005
R7600 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 17.4005
R7601 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 17.2391
R7602 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 9.52217
R7603 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 9.52217
R7604 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 6.39571
R7605 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 5.30824
R7606 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 4.94887
R7607 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 1.06691
R7608 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 890.727
R7609 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 742.783
R7610 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 641.061
R7611 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7612 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 547.874
R7613 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7614 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 427.875
R7615 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7616 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7617 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7618 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7619 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R7620 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 31.0962
R7621 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R7622 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7623 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 8.91506
R7624 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7625 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7626 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7627 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7628 uo_out[5].n0 uo_out[5].t4 734.539
R7629 uo_out[5].n0 uo_out[5].t5 233.26
R7630 uo_out[5].n2 uo_out[5].n0 162.335
R7631 uo_out[5].n2 uo_out[5].n1 75.5733
R7632 uo_out[5].n4 uo_out[5].n3 66.3172
R7633 uo_out[5].n5 uo_out[5] 19.2682
R7634 uo_out[5].n3 uo_out[5].t1 17.4005
R7635 uo_out[5].n3 uo_out[5].t2 17.4005
R7636 uo_out[5].n1 uo_out[5].t3 9.52217
R7637 uo_out[5].n1 uo_out[5].t0 9.52217
R7638 uo_out[5].n5 uo_out[5].n4 5.02496
R7639 uo_out[5].n4 uo_out[5].n2 0.438
R7640 uo_out[5] uo_out[5].n5 0.063
R7641 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 552.84
R7642 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 552.84
R7643 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 552.84
R7644 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 552.84
R7645 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 539.841
R7646 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 539.841
R7647 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 539.841
R7648 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 539.841
R7649 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 215.293
R7650 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 215.293
R7651 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 215.293
R7652 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 215.293
R7653 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 166.468
R7654 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 166.149
R7655 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 165.8
R7656 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 165.8
R7657 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 85.1574
R7658 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 83.8097
R7659 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 83.8097
R7660 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 83.7172
R7661 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 74.288
R7662 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 67.7574
R7663 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 36.1505
R7664 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 36.1505
R7665 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 34.5438
R7666 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 34.5438
R7667 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 17.4005
R7668 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 17.4005
R7669 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 16.09
R7670 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 11.8364
R7671 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 9.52217
R7672 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 9.52217
R7673 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 5.96628
R7674 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 5.83219
R7675 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 5.74235
R7676 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 5.49235
R7677 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 1.44072
R7678 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 1.32081
R7679 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 0.285656
R7680 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 628.097
R7681 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 622.766
R7682 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 523.774
R7683 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 304.647
R7684 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 304.647
R7685 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 202.44
R7686 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 169.062
R7687 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 166.237
R7688 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 84.7557
R7689 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 84.1197
R7690 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 12.6535
R7691 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 5.48979
R7692 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 4.5005
R7693 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 1.09595
R7694 ui_in[5].n0 ui_in[5].t7 628.097
R7695 ui_in[5].n1 ui_in[5].t3 622.766
R7696 ui_in[5].n5 ui_in[5].t0 543.053
R7697 ui_in[5].n0 ui_in[5].t5 523.774
R7698 ui_in[5].n2 ui_in[5].t6 304.647
R7699 ui_in[5].n2 ui_in[5].t2 304.647
R7700 ui_in[5].n5 ui_in[5].t1 221.72
R7701 ui_in[5].n6 ui_in[5].n5 220.327
R7702 ui_in[5].n2 ui_in[5].t4 202.44
R7703 ui_in[5] ui_in[5].n2 169.071
R7704 ui_in[5] ui_in[5].n1 166.244
R7705 ui_in[5].n4 ui_in[5] 30.5822
R7706 ui_in[5].n4 ui_in[5].n3 3.0755
R7707 ui_in[5].n3 ui_in[5] 1.24128
R7708 ui_in[5].n1 ui_in[5].n0 1.09595
R7709 ui_in[5].n3 ui_in[5] 0.402286
R7710 ui_in[5].n6 ui_in[5] 0.063
R7711 ui_in[5] ui_in[5].n6 0.0505
R7712 ui_in[5] ui_in[5].n4 0.0147857
R7713 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 539.841
R7714 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 539.841
R7715 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 539.841
R7716 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 539.841
R7717 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 215.293
R7718 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 215.293
R7719 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 215.293
R7720 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 215.293
R7721 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 166.144
R7722 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 165.8
R7723 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 85.2499
R7724 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 85.2499
R7725 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 83.7172
R7726 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 83.7172
R7727 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 75.7282
R7728 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 66.3172
R7729 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 36.1505
R7730 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 36.1505
R7731 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 34.5438
R7732 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 34.5438
R7733 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 17.4005
R7734 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 17.4005
R7735 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 9.52217
R7736 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 9.52217
R7737 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 6.39571
R7738 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 5.30824
R7739 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 4.94887
R7740 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 1.06691
R7741 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 0.160656
R7742 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 539.841
R7743 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 539.841
R7744 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 539.841
R7745 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 539.841
R7746 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 215.293
R7747 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 215.293
R7748 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 215.293
R7749 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 215.293
R7750 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 166.149
R7751 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 165.8
R7752 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 85.1574
R7753 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 85.1574
R7754 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 83.8097
R7755 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 83.8097
R7756 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 74.288
R7757 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 67.7574
R7758 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 36.1505
R7759 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 36.1505
R7760 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 34.5438
R7761 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 34.5438
R7762 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 17.4005
R7763 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 17.4005
R7764 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 11.8364
R7765 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 9.52217
R7766 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 9.52217
R7767 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 5.83219
R7768 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 5.74235
R7769 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 5.49235
R7770 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 1.32081
R7771 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 0.285656
R7772 a_10958_27928.n2 a_10958_27928.t3 31.9657
R7773 a_10958_27928.n2 a_10958_27928.n1 25.8125
R7774 a_10958_27928.n4 a_10958_27928.n3 25.8125
R7775 a_10958_27928.n6 a_10958_27928.n5 25.8125
R7776 a_10958_27928.n9 a_10958_27928.n0 25.7038
R7777 a_10958_27928.n10 a_10958_27928.n9 25.3505
R7778 a_10958_27928.n8 a_10958_27928.n7 24.288
R7779 a_10958_27928.n7 a_10958_27928.t6 5.8005
R7780 a_10958_27928.n7 a_10958_27928.t10 5.8005
R7781 a_10958_27928.n1 a_10958_27928.t11 5.8005
R7782 a_10958_27928.n1 a_10958_27928.t0 5.8005
R7783 a_10958_27928.n3 a_10958_27928.t2 5.8005
R7784 a_10958_27928.n3 a_10958_27928.t9 5.8005
R7785 a_10958_27928.n5 a_10958_27928.t12 5.8005
R7786 a_10958_27928.n5 a_10958_27928.t1 5.8005
R7787 a_10958_27928.n0 a_10958_27928.t4 5.8005
R7788 a_10958_27928.n0 a_10958_27928.t7 5.8005
R7789 a_10958_27928.t8 a_10958_27928.n10 5.8005
R7790 a_10958_27928.n10 a_10958_27928.t5 5.8005
R7791 a_10958_27928.n8 a_10958_27928.n6 1.87822
R7792 a_10958_27928.n9 a_10958_27928.n8 1.41626
R7793 a_10958_27928.n4 a_10958_27928.n2 0.353761
R7794 a_10958_27928.n6 a_10958_27928.n4 0.353761
R7795 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 879.481
R7796 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7797 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 641.061
R7798 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 623.388
R7799 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 547.874
R7800 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 431.807
R7801 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 427.875
R7802 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7803 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7804 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7805 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7806 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7807 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 31.2972
R7808 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 11.1806
R7809 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7810 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R7811 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R7812 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7813 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 628.097
R7814 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 622.766
R7815 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 523.774
R7816 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 304.647
R7817 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 304.647
R7818 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 202.44
R7819 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 169.062
R7820 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 166.237
R7821 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 84.7557
R7822 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 84.1197
R7823 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R7824 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 5.48979
R7825 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en 4.5005
R7826 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 1.09595
R7827 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 784.053
R7828 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 784.053
R7829 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 784.053
R7830 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 784.053
R7831 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 539.841
R7832 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 539.841
R7833 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 539.841
R7834 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 539.841
R7835 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 215.293
R7836 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 215.293
R7837 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 215.293
R7838 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 215.293
R7839 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 168.659
R7840 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 167.992
R7841 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 166.144
R7842 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 165.8
R7843 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 85.2499
R7844 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 85.2499
R7845 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 83.7172
R7846 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 83.7172
R7847 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 75.7282
R7848 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 66.3172
R7849 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 36.1505
R7850 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 36.1505
R7851 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 34.5438
R7852 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 34.5438
R7853 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 17.4005
R7854 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 17.4005
R7855 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 17.2391
R7856 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 9.52217
R7857 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 9.52217
R7858 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 6.39571
R7859 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 5.30824
R7860 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 4.94887
R7861 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 1.06691
R7862 a_10108_30826.n2 a_10108_30826.n1 34.9195
R7863 a_10108_30826.n3 a_10108_30826.n2 25.5407
R7864 a_10108_30826.n2 a_10108_30826.n0 25.2907
R7865 a_10108_30826.n1 a_10108_30826.t1 5.8005
R7866 a_10108_30826.n1 a_10108_30826.t2 5.8005
R7867 a_10108_30826.n0 a_10108_30826.t0 5.8005
R7868 a_10108_30826.n0 a_10108_30826.t3 5.8005
R7869 a_10108_30826.t4 a_10108_30826.n3 5.8005
R7870 a_10108_30826.n3 a_10108_30826.t5 5.8005
R7871 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 784.053
R7872 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 784.053
R7873 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 784.053
R7874 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 784.053
R7875 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 539.841
R7876 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 539.841
R7877 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 539.841
R7878 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 539.841
R7879 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 215.293
R7880 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 215.293
R7881 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 215.293
R7882 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 215.293
R7883 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 168.659
R7884 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 167.992
R7885 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 166.144
R7886 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 165.8
R7887 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 85.2499
R7888 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 85.2499
R7889 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 83.7172
R7890 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 83.7172
R7891 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 75.7282
R7892 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 66.3172
R7893 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 36.1505
R7894 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 36.1505
R7895 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 34.5438
R7896 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 34.5438
R7897 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 17.4005
R7898 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 17.4005
R7899 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 17.2391
R7900 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 9.52217
R7901 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 9.52217
R7902 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 6.39571
R7903 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 5.30824
R7904 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 4.94887
R7905 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 1.06691
R7906 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 539.841
R7907 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 539.841
R7908 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 539.841
R7909 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 539.841
R7910 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 215.293
R7911 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 215.293
R7912 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 215.293
R7913 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 215.293
R7914 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 166.149
R7915 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 165.8
R7916 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 85.1574
R7917 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 85.1574
R7918 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 83.8097
R7919 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 83.8097
R7920 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 74.288
R7921 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 67.7574
R7922 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 36.1505
R7923 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 36.1505
R7924 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 34.5438
R7925 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 34.5438
R7926 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 17.4005
R7927 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 17.4005
R7928 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 11.8364
R7929 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 9.52217
R7930 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 9.52217
R7931 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 5.83219
R7932 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 5.74235
R7933 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 5.49235
R7934 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 1.32081
R7935 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 0.285656
R7936 uo_out[0].n0 uo_out[0].t5 734.539
R7937 uo_out[0].n0 uo_out[0].t4 233.26
R7938 uo_out[0].n2 uo_out[0].n0 162.335
R7939 uo_out[0].n2 uo_out[0].n1 75.5733
R7940 uo_out[0].n4 uo_out[0].n3 66.3172
R7941 uo_out[0].n5 uo_out[0] 33.5966
R7942 uo_out[0].n3 uo_out[0].t2 17.4005
R7943 uo_out[0].n3 uo_out[0].t0 17.4005
R7944 uo_out[0].n1 uo_out[0].t1 9.52217
R7945 uo_out[0].n1 uo_out[0].t3 9.52217
R7946 uo_out[0].n5 uo_out[0].n4 5.02496
R7947 uo_out[0].n4 uo_out[0].n2 0.438
R7948 uo_out[0] uo_out[0].n5 0.063
R7949 a_10958_25646.n1 a_10958_25646.t4 31.9657
R7950 a_10958_25646.n1 a_10958_25646.n0 25.8125
R7951 a_10958_25646.n3 a_10958_25646.n2 25.8125
R7952 a_10958_25646.n5 a_10958_25646.n4 25.8125
R7953 a_10958_25646.n8 a_10958_25646.n6 25.7038
R7954 a_10958_25646.n8 a_10958_25646.n7 25.3505
R7955 a_10958_25646.n10 a_10958_25646.n9 24.288
R7956 a_10958_25646.n6 a_10958_25646.t9 5.8005
R7957 a_10958_25646.n6 a_10958_25646.t10 5.8005
R7958 a_10958_25646.n7 a_10958_25646.t7 5.8005
R7959 a_10958_25646.n7 a_10958_25646.t8 5.8005
R7960 a_10958_25646.n0 a_10958_25646.t2 5.8005
R7961 a_10958_25646.n0 a_10958_25646.t5 5.8005
R7962 a_10958_25646.n2 a_10958_25646.t12 5.8005
R7963 a_10958_25646.n2 a_10958_25646.t1 5.8005
R7964 a_10958_25646.n4 a_10958_25646.t0 5.8005
R7965 a_10958_25646.n4 a_10958_25646.t6 5.8005
R7966 a_10958_25646.t11 a_10958_25646.n10 5.8005
R7967 a_10958_25646.n10 a_10958_25646.t3 5.8005
R7968 a_10958_25646.n9 a_10958_25646.n5 1.87822
R7969 a_10958_25646.n9 a_10958_25646.n8 1.41626
R7970 a_10958_25646.n3 a_10958_25646.n1 0.353761
R7971 a_10958_25646.n5 a_10958_25646.n3 0.353761
R7972 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 890.727
R7973 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 742.783
R7974 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 641.061
R7975 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 623.388
R7976 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 547.874
R7977 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 431.807
R7978 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 427.875
R7979 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7980 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7981 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7982 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7983 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 31.2103
R7984 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 31.0962
R7985 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7986 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R7987 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 8.91506
R7988 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7989 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7990 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7991 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7992 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 879.481
R7993 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 742.783
R7994 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 641.061
R7995 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 623.388
R7996 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 547.874
R7997 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 431.807
R7998 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 427.875
R7999 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 333.161
R8000 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 208.668
R8001 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 168.077
R8002 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 75.5951
R8003 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R8004 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R8005 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 11.1806
R8006 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 10.4291
R8007 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8008 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R8009 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 0.740618
R8010 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 0.228761
R8011 uo_out[3].n0 uo_out[3].t4 734.539
R8012 uo_out[3].n0 uo_out[3].t5 233.26
R8013 uo_out[3].n2 uo_out[3].n0 162.335
R8014 uo_out[3].n2 uo_out[3].n1 75.5733
R8015 uo_out[3].n4 uo_out[3].n3 66.3172
R8016 uo_out[3].n5 uo_out[3] 24.9996
R8017 uo_out[3].n3 uo_out[3].t0 17.4005
R8018 uo_out[3].n3 uo_out[3].t2 17.4005
R8019 uo_out[3].n1 uo_out[3].t3 9.52217
R8020 uo_out[3].n1 uo_out[3].t1 9.52217
R8021 uo_out[3].n5 uo_out[3].n4 5.02496
R8022 uo_out[3].n4 uo_out[3].n2 0.438
R8023 uo_out[3] uo_out[3].n5 0.063
R8024 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 628.097
R8025 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 622.766
R8026 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 523.774
R8027 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 304.647
R8028 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 304.647
R8029 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 202.44
R8030 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 169.062
R8031 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 166.237
R8032 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R8033 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R8034 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R8035 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 5.48979
R8036 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 4.5005
R8037 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 1.09595
R8038 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 539.841
R8039 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 539.841
R8040 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 539.841
R8041 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 539.841
R8042 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 215.293
R8043 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 215.293
R8044 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 215.293
R8045 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 215.293
R8046 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 166.144
R8047 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 165.8
R8048 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 85.2499
R8049 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 85.2499
R8050 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 83.7172
R8051 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 83.7172
R8052 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 75.7282
R8053 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 66.3172
R8054 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 36.1505
R8055 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 36.1505
R8056 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 34.5438
R8057 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 34.5438
R8058 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 17.4005
R8059 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 17.4005
R8060 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 9.52217
R8061 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 9.52217
R8062 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 6.39571
R8063 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 5.30824
R8064 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 4.94887
R8065 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 1.41456
R8066 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 539.841
R8067 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 539.841
R8068 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 539.841
R8069 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 539.841
R8070 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 215.293
R8071 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 215.293
R8072 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 215.293
R8073 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 215.293
R8074 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 166.149
R8075 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 165.8
R8076 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 85.1574
R8077 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 85.1574
R8078 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 83.8097
R8079 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 83.8097
R8080 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 74.288
R8081 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 67.7574
R8082 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 36.1505
R8083 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 36.1505
R8084 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 34.5438
R8085 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 34.5438
R8086 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 17.4005
R8087 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 17.4005
R8088 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 11.8364
R8089 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 9.52217
R8090 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 9.52217
R8091 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 5.83219
R8092 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 5.74235
R8093 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 5.49235
R8094 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 1.32081
R8095 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 0.285656
R8096 a_10958_32492.n1 a_10958_32492.t11 31.9657
R8097 a_10958_32492.n1 a_10958_32492.n0 25.8125
R8098 a_10958_32492.n3 a_10958_32492.n2 25.8125
R8099 a_10958_32492.n5 a_10958_32492.n4 25.8125
R8100 a_10958_32492.n10 a_10958_32492.n9 25.7038
R8101 a_10958_32492.n9 a_10958_32492.n8 25.3505
R8102 a_10958_32492.n7 a_10958_32492.n6 24.288
R8103 a_10958_32492.n6 a_10958_32492.t8 5.8005
R8104 a_10958_32492.n6 a_10958_32492.t0 5.8005
R8105 a_10958_32492.n0 a_10958_32492.t1 5.8005
R8106 a_10958_32492.n0 a_10958_32492.t12 5.8005
R8107 a_10958_32492.n2 a_10958_32492.t10 5.8005
R8108 a_10958_32492.n2 a_10958_32492.t4 5.8005
R8109 a_10958_32492.n4 a_10958_32492.t3 5.8005
R8110 a_10958_32492.n4 a_10958_32492.t2 5.8005
R8111 a_10958_32492.n8 a_10958_32492.t6 5.8005
R8112 a_10958_32492.n8 a_10958_32492.t7 5.8005
R8113 a_10958_32492.t9 a_10958_32492.n10 5.8005
R8114 a_10958_32492.n10 a_10958_32492.t5 5.8005
R8115 a_10958_32492.n7 a_10958_32492.n5 1.87822
R8116 a_10958_32492.n9 a_10958_32492.n7 1.41626
R8117 a_10958_32492.n3 a_10958_32492.n1 0.353761
R8118 a_10958_32492.n5 a_10958_32492.n3 0.353761
R8119 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 552.84
R8120 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 552.84
R8121 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 552.84
R8122 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 552.84
R8123 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 539.841
R8124 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 539.841
R8125 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 539.841
R8126 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 539.841
R8127 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 215.293
R8128 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 215.293
R8129 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 215.293
R8130 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 215.293
R8131 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 166.468
R8132 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 166.149
R8133 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 165.8
R8134 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 165.8
R8135 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 85.1574
R8136 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 83.8097
R8137 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 83.8097
R8138 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 83.7172
R8139 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 74.288
R8140 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 67.7574
R8141 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 36.1505
R8142 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 36.1505
R8143 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 34.5438
R8144 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 34.5438
R8145 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 17.4005
R8146 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 17.4005
R8147 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 16.09
R8148 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 11.8364
R8149 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 9.52217
R8150 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 9.52217
R8151 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 5.96628
R8152 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 5.83219
R8153 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 5.74235
R8154 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 5.49235
R8155 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 1.44072
R8156 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 1.32081
R8157 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 539.841
R8158 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 539.841
R8159 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 539.841
R8160 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 539.841
R8161 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 215.293
R8162 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 215.293
R8163 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 215.293
R8164 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 215.293
R8165 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 166.149
R8166 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 165.8
R8167 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 85.1574
R8168 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 85.1574
R8169 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 83.8097
R8170 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 83.8097
R8171 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 74.288
R8172 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 67.7574
R8173 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 36.1505
R8174 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 36.1505
R8175 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 34.5438
R8176 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 34.5438
R8177 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 17.4005
R8178 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 17.4005
R8179 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 11.8364
R8180 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 9.52217
R8181 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 9.52217
R8182 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 5.83219
R8183 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 5.74235
R8184 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 5.49235
R8185 tdc_0.diff_gen_0.delay_unit_2_1.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 1.32081
R8186 tdc_0.diff_gen_0.delay_unit_2_1.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 0.285656
R8187 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 784.053
R8188 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 784.053
R8189 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 784.053
R8190 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 784.053
R8191 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 539.841
R8192 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 539.841
R8193 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 539.841
R8194 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 539.841
R8195 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 215.293
R8196 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 215.293
R8197 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 215.293
R8198 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 215.293
R8199 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 168.659
R8200 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 167.992
R8201 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 166.144
R8202 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 165.8
R8203 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 85.2499
R8204 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 85.2499
R8205 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 83.7172
R8206 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 83.7172
R8207 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 75.7282
R8208 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 66.3172
R8209 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 36.1505
R8210 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 36.1505
R8211 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 34.5438
R8212 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 34.5438
R8213 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 17.4005
R8214 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 17.4005
R8215 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 17.2391
R8216 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 9.52217
R8217 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 9.52217
R8218 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 6.39571
R8219 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 5.30824
R8220 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 4.94887
R8221 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 1.06691
R8222 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 879.481
R8223 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 742.783
R8224 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 641.061
R8225 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 623.388
R8226 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 547.874
R8227 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 431.807
R8228 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 427.875
R8229 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 333.161
R8230 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 208.668
R8231 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 168.077
R8232 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R8233 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R8234 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R8235 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 11.1806
R8236 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R8237 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8238 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R8239 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R8240 variable_delay_short_0.variable_delay_unit_5.in.n0 variable_delay_short_0.variable_delay_unit_5.in.t5 607.409
R8241 variable_delay_short_0.variable_delay_unit_5.in.n2 variable_delay_short_0.variable_delay_unit_5.in.t2 543.053
R8242 variable_delay_short_0.variable_delay_unit_5.in.n0 variable_delay_short_0.variable_delay_unit_5.in.t4 321.423
R8243 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n2 221.778
R8244 variable_delay_short_0.variable_delay_unit_5.in.n2 variable_delay_short_0.variable_delay_unit_5.in.t3 221.72
R8245 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n0 161.72
R8246 variable_delay_short_0.variable_delay_unit_5.in.n1 variable_delay_short_0.variable_delay_unit_5.in.t1 84.7227
R8247 variable_delay_short_0.variable_delay_unit_5.in.n1 variable_delay_short_0.variable_delay_unit_5.in.t0 84.0867
R8248 variable_delay_short_0.variable_delay_unit_5.in.n3 variable_delay_short_0.variable_delay_unit_5.in 20.0791
R8249 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n3 0.851271
R8250 variable_delay_short_0.variable_delay_unit_5.in.n3 variable_delay_short_0.variable_delay_unit_5.in.n1 0.465495
R8251 variable_delay_short_0.variable_delay_unit_5.forward.n0 variable_delay_short_0.variable_delay_unit_5.forward.t3 607.409
R8252 variable_delay_short_0.variable_delay_unit_5.forward.n0 variable_delay_short_0.variable_delay_unit_5.forward.t2 321.423
R8253 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.forward.n0 161.72
R8254 variable_delay_short_0.variable_delay_unit_5.forward.n1 variable_delay_short_0.variable_delay_unit_5.forward.t1 84.7227
R8255 variable_delay_short_0.variable_delay_unit_5.forward.n1 variable_delay_short_0.variable_delay_unit_5.forward.t0 84.0867
R8256 variable_delay_short_0.variable_delay_unit_5.forward.n2 variable_delay_short_0.variable_delay_unit_5.forward 19.7898
R8257 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.forward.n2 0.851271
R8258 variable_delay_short_0.variable_delay_unit_5.forward.n2 variable_delay_short_0.variable_delay_unit_5.forward.n1 0.465495
R8259 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 552.84
R8260 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 552.84
R8261 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 552.84
R8262 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 552.84
R8263 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 539.841
R8264 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 539.841
R8265 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 539.841
R8266 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 539.841
R8267 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 215.293
R8268 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 215.293
R8269 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 215.293
R8270 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 215.293
R8271 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 166.468
R8272 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 166.149
R8273 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 165.8
R8274 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 165.8
R8275 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 85.1574
R8276 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 83.8097
R8277 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 83.8097
R8278 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 83.7172
R8279 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 74.288
R8280 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 67.7574
R8281 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 36.1505
R8282 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 36.1505
R8283 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 34.5438
R8284 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 34.5438
R8285 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 17.4005
R8286 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 17.4005
R8287 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 16.09
R8288 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 11.8364
R8289 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 9.52217
R8290 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 9.52217
R8291 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 5.96628
R8292 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 5.83219
R8293 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 5.74235
R8294 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 5.49235
R8295 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 1.44072
R8296 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 1.32081
R8297 a_10958_30210.n2 a_10958_30210.t12 31.9657
R8298 a_10958_30210.n2 a_10958_30210.n1 25.8125
R8299 a_10958_30210.n4 a_10958_30210.n3 25.8125
R8300 a_10958_30210.n6 a_10958_30210.n5 25.8125
R8301 a_10958_30210.n9 a_10958_30210.n0 25.7038
R8302 a_10958_30210.n10 a_10958_30210.n9 25.3505
R8303 a_10958_30210.n8 a_10958_30210.n7 24.288
R8304 a_10958_30210.n7 a_10958_30210.t1 5.8005
R8305 a_10958_30210.n7 a_10958_30210.t6 5.8005
R8306 a_10958_30210.n1 a_10958_30210.t5 5.8005
R8307 a_10958_30210.n1 a_10958_30210.t9 5.8005
R8308 a_10958_30210.n3 a_10958_30210.t11 5.8005
R8309 a_10958_30210.n3 a_10958_30210.t7 5.8005
R8310 a_10958_30210.n5 a_10958_30210.t8 5.8005
R8311 a_10958_30210.n5 a_10958_30210.t10 5.8005
R8312 a_10958_30210.n0 a_10958_30210.t0 5.8005
R8313 a_10958_30210.n0 a_10958_30210.t2 5.8005
R8314 a_10958_30210.n10 a_10958_30210.t3 5.8005
R8315 a_10958_30210.t4 a_10958_30210.n10 5.8005
R8316 a_10958_30210.n8 a_10958_30210.n6 1.87822
R8317 a_10958_30210.n9 a_10958_30210.n8 1.41626
R8318 a_10958_30210.n4 a_10958_30210.n2 0.353761
R8319 a_10958_30210.n6 a_10958_30210.n4 0.353761
R8320 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 784.053
R8321 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 784.053
R8322 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 784.053
R8323 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 784.053
R8324 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 539.841
R8325 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 539.841
R8326 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 539.841
R8327 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 539.841
R8328 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 215.293
R8329 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 215.293
R8330 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 215.293
R8331 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 215.293
R8332 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 168.659
R8333 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 167.992
R8334 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 166.144
R8335 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 165.8
R8336 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 85.2499
R8337 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 85.2499
R8338 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 83.7172
R8339 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 83.7172
R8340 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 75.7282
R8341 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 66.3172
R8342 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 36.1505
R8343 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 36.1505
R8344 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 34.5438
R8345 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 34.5438
R8346 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 17.4005
R8347 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 17.4005
R8348 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 17.2391
R8349 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 9.52217
R8350 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 9.52217
R8351 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 6.39571
R8352 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 5.30824
R8353 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 4.94887
R8354 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 1.06691
R8355 a_10108_23980.n2 a_10108_23980.n1 34.9195
R8356 a_10108_23980.n2 a_10108_23980.n0 25.5407
R8357 a_10108_23980.n3 a_10108_23980.n2 25.2907
R8358 a_10108_23980.n1 a_10108_23980.t3 5.8005
R8359 a_10108_23980.n1 a_10108_23980.t5 5.8005
R8360 a_10108_23980.n0 a_10108_23980.t0 5.8005
R8361 a_10108_23980.n0 a_10108_23980.t1 5.8005
R8362 a_10108_23980.n3 a_10108_23980.t2 5.8005
R8363 a_10108_23980.t4 a_10108_23980.n3 5.8005
R8364 variable_delay_short_0.variable_delay_unit_3.in.n0 variable_delay_short_0.variable_delay_unit_3.in.t5 607.409
R8365 variable_delay_short_0.variable_delay_unit_3.in.n2 variable_delay_short_0.variable_delay_unit_3.in.t2 543.053
R8366 variable_delay_short_0.variable_delay_unit_3.in.n0 variable_delay_short_0.variable_delay_unit_3.in.t4 321.423
R8367 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n2 221.778
R8368 variable_delay_short_0.variable_delay_unit_3.in.n2 variable_delay_short_0.variable_delay_unit_3.in.t3 221.72
R8369 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n0 161.72
R8370 variable_delay_short_0.variable_delay_unit_3.in.n1 variable_delay_short_0.variable_delay_unit_3.in.t1 84.7227
R8371 variable_delay_short_0.variable_delay_unit_3.in.n1 variable_delay_short_0.variable_delay_unit_3.in.t0 84.0867
R8372 variable_delay_short_0.variable_delay_unit_3.in.n3 variable_delay_short_0.variable_delay_unit_3.in 20.0791
R8373 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n3 0.851271
R8374 variable_delay_short_0.variable_delay_unit_3.in.n3 variable_delay_short_0.variable_delay_unit_3.in.n1 0.465495
R8375 variable_delay_short_0.variable_delay_unit_4.in.n0 variable_delay_short_0.variable_delay_unit_4.in.t5 607.409
R8376 variable_delay_short_0.variable_delay_unit_4.in.n2 variable_delay_short_0.variable_delay_unit_4.in.t2 543.053
R8377 variable_delay_short_0.variable_delay_unit_4.in.n0 variable_delay_short_0.variable_delay_unit_4.in.t4 321.423
R8378 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n2 221.778
R8379 variable_delay_short_0.variable_delay_unit_4.in.n2 variable_delay_short_0.variable_delay_unit_4.in.t3 221.72
R8380 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n0 161.72
R8381 variable_delay_short_0.variable_delay_unit_4.in.n1 variable_delay_short_0.variable_delay_unit_4.in.t1 84.7227
R8382 variable_delay_short_0.variable_delay_unit_4.in.n1 variable_delay_short_0.variable_delay_unit_4.in.t0 84.0867
R8383 variable_delay_short_0.variable_delay_unit_4.in.n3 variable_delay_short_0.variable_delay_unit_4.in 20.0791
R8384 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n3 0.851271
R8385 variable_delay_short_0.variable_delay_unit_4.in.n3 variable_delay_short_0.variable_delay_unit_4.in.n1 0.465495
R8386 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 552.84
R8387 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 552.84
R8388 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 552.84
R8389 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 552.84
R8390 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 539.841
R8391 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 539.841
R8392 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 539.841
R8393 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 539.841
R8394 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 215.293
R8395 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 215.293
R8396 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 215.293
R8397 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 215.293
R8398 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 166.468
R8399 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 166.149
R8400 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 165.8
R8401 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 165.8
R8402 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 85.1574
R8403 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 83.8097
R8404 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 83.8097
R8405 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 83.7172
R8406 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 74.288
R8407 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 67.7574
R8408 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 36.1505
R8409 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 36.1505
R8410 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 34.5438
R8411 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 34.5438
R8412 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 17.4005
R8413 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 17.4005
R8414 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 16.09
R8415 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 11.8364
R8416 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 9.52217
R8417 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 9.52217
R8418 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 5.96628
R8419 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 5.83219
R8420 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 5.74235
R8421 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 5.49235
R8422 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 1.44072
R8423 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 1.32081
R8424 uo_out[4].n0 uo_out[4].t5 734.539
R8425 uo_out[4].n0 uo_out[4].t4 233.26
R8426 uo_out[4].n2 uo_out[4].n0 162.335
R8427 uo_out[4].n2 uo_out[4].n1 75.5733
R8428 uo_out[4].n4 uo_out[4].n3 66.3172
R8429 uo_out[4].n5 uo_out[4] 22.1339
R8430 uo_out[4].n3 uo_out[4].t3 17.4005
R8431 uo_out[4].n3 uo_out[4].t0 17.4005
R8432 uo_out[4].n1 uo_out[4].t1 9.52217
R8433 uo_out[4].n1 uo_out[4].t2 9.52217
R8434 uo_out[4].n5 uo_out[4].n4 5.02496
R8435 uo_out[4].n4 uo_out[4].n2 0.438
R8436 uo_out[4] uo_out[4].n5 0.063
R8437 ui_in[4].n1 ui_in[4].t2 628.097
R8438 ui_in[4].n2 ui_in[4].t6 622.766
R8439 ui_in[4].n0 ui_in[4].t3 543.053
R8440 ui_in[4].n1 ui_in[4].t0 523.774
R8441 ui_in[4].n3 ui_in[4].t1 304.647
R8442 ui_in[4].n3 ui_in[4].t4 304.647
R8443 ui_in[4].n0 ui_in[4].t5 221.72
R8444 ui_in[4].n6 ui_in[4].n0 220.327
R8445 ui_in[4].n3 ui_in[4].t7 202.44
R8446 ui_in[4] ui_in[4].n3 169.071
R8447 ui_in[4] ui_in[4].n2 166.244
R8448 ui_in[4].n5 ui_in[4] 27.1791
R8449 ui_in[4].n5 ui_in[4].n4 2.98979
R8450 ui_in[4].n4 ui_in[4] 1.24128
R8451 ui_in[4].n2 ui_in[4].n1 1.09595
R8452 ui_in[4].n4 ui_in[4] 0.402286
R8453 ui_in[4].n6 ui_in[4].n5 0.1505
R8454 ui_in[4].n6 ui_in[4] 0.063
R8455 ui_in[4] ui_in[4].n6 0.0219286
R8456 uo_out[7].n0 uo_out[7].t5 734.539
R8457 uo_out[7].n0 uo_out[7].t4 233.26
R8458 uo_out[7].n2 uo_out[7].n0 162.335
R8459 uo_out[7].n2 uo_out[7].n1 75.5733
R8460 uo_out[7].n4 uo_out[7].n3 66.3172
R8461 uo_out[7].n3 uo_out[7].t1 17.4005
R8462 uo_out[7].n3 uo_out[7].t2 17.4005
R8463 uo_out[7].n5 uo_out[7] 13.5368
R8464 uo_out[7].n1 uo_out[7].t3 9.52217
R8465 uo_out[7].n1 uo_out[7].t0 9.52217
R8466 uo_out[7].n5 uo_out[7].n4 5.02496
R8467 uo_out[7].n4 uo_out[7].n2 0.438
R8468 uo_out[7] uo_out[7].n5 0.063
R8469 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 552.84
R8470 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 552.84
R8471 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 552.84
R8472 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 552.84
R8473 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 539.841
R8474 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 539.841
R8475 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 539.841
R8476 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 539.841
R8477 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 215.293
R8478 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 215.293
R8479 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 215.293
R8480 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 215.293
R8481 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 166.468
R8482 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 166.149
R8483 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 165.8
R8484 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 165.8
R8485 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 85.1574
R8486 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 83.8097
R8487 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 83.8097
R8488 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 83.7172
R8489 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 74.288
R8490 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 67.7574
R8491 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 36.1505
R8492 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 36.1505
R8493 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 34.5438
R8494 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 34.5438
R8495 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 17.4005
R8496 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 17.4005
R8497 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 16.09
R8498 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 11.8364
R8499 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 9.52217
R8500 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 9.52217
R8501 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 5.96628
R8502 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 5.83219
R8503 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 5.74235
R8504 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 5.49235
R8505 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 1.44072
R8506 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 1.32081
R8507 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 0.285656
R8508 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 539.841
R8509 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 539.841
R8510 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 539.841
R8511 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 539.841
R8512 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 215.293
R8513 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 215.293
R8514 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 215.293
R8515 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 215.293
R8516 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 166.144
R8517 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 165.8
R8518 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 85.2499
R8519 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 85.2499
R8520 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 83.7172
R8521 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 83.7172
R8522 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 75.7282
R8523 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 66.3172
R8524 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 36.1505
R8525 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 36.1505
R8526 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 34.5438
R8527 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 34.5438
R8528 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 17.4005
R8529 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 17.4005
R8530 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 9.52217
R8531 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 9.52217
R8532 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 6.39571
R8533 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 5.30824
R8534 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 4.94887
R8535 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 1.06691
R8536 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 0.160656
R8537 tdc_0.vernier_delay_line_0.start_pos.n1 tdc_0.vernier_delay_line_0.start_pos.t8 539.841
R8538 tdc_0.vernier_delay_line_0.start_pos.n0 tdc_0.vernier_delay_line_0.start_pos.t11 539.841
R8539 tdc_0.vernier_delay_line_0.start_pos.n4 tdc_0.vernier_delay_line_0.start_pos.t12 539.841
R8540 tdc_0.vernier_delay_line_0.start_pos.n3 tdc_0.vernier_delay_line_0.start_pos.t14 539.841
R8541 tdc_0.vernier_delay_line_0.start_pos.n1 tdc_0.vernier_delay_line_0.start_pos.t15 215.293
R8542 tdc_0.vernier_delay_line_0.start_pos.n0 tdc_0.vernier_delay_line_0.start_pos.t9 215.293
R8543 tdc_0.vernier_delay_line_0.start_pos.n4 tdc_0.vernier_delay_line_0.start_pos.t10 215.293
R8544 tdc_0.vernier_delay_line_0.start_pos.n3 tdc_0.vernier_delay_line_0.start_pos.t13 215.293
R8545 tdc_0.vernier_delay_line_0.start_pos.n6 tdc_0.vernier_delay_line_0.start_pos.n2 166.149
R8546 tdc_0.vernier_delay_line_0.start_pos.n6 tdc_0.vernier_delay_line_0.start_pos.n5 165.8
R8547 tdc_0.vernier_delay_line_0.start_pos.n12 tdc_0.vernier_delay_line_0.start_pos.t0 85.1574
R8548 tdc_0.vernier_delay_line_0.start_pos.n7 tdc_0.vernier_delay_line_0.start_pos.t6 85.1574
R8549 tdc_0.vernier_delay_line_0.start_pos.n7 tdc_0.vernier_delay_line_0.start_pos.t7 83.8097
R8550 tdc_0.vernier_delay_line_0.start_pos.n12 tdc_0.vernier_delay_line_0.start_pos.t5 83.8097
R8551 tdc_0.vernier_delay_line_0.start_pos.n11 tdc_0.vernier_delay_line_0.start_pos.n10 74.288
R8552 tdc_0.vernier_delay_line_0.start_pos.n11 tdc_0.vernier_delay_line_0.start_pos.n9 67.7574
R8553 tdc_0.vernier_delay_line_0.start_pos.n2 tdc_0.vernier_delay_line_0.start_pos.n1 36.1505
R8554 tdc_0.vernier_delay_line_0.start_pos.n5 tdc_0.vernier_delay_line_0.start_pos.n3 36.1505
R8555 tdc_0.vernier_delay_line_0.start_pos.n2 tdc_0.vernier_delay_line_0.start_pos.n0 34.5438
R8556 tdc_0.vernier_delay_line_0.start_pos.n5 tdc_0.vernier_delay_line_0.start_pos.n4 34.5438
R8557 tdc_0.vernier_delay_line_0.start_pos.n9 tdc_0.vernier_delay_line_0.start_pos.t1 17.4005
R8558 tdc_0.vernier_delay_line_0.start_pos.n9 tdc_0.vernier_delay_line_0.start_pos.t2 17.4005
R8559 tdc_0.vernier_delay_line_0.start_pos.n8 tdc_0.vernier_delay_line_0.start_pos.n6 11.8364
R8560 tdc_0.vernier_delay_line_0.start_pos.n10 tdc_0.vernier_delay_line_0.start_pos.t3 9.52217
R8561 tdc_0.vernier_delay_line_0.start_pos.n10 tdc_0.vernier_delay_line_0.start_pos.t4 9.52217
R8562 tdc_0.vernier_delay_line_0.start_pos.n13 tdc_0.vernier_delay_line_0.start_pos.n11 5.83219
R8563 tdc_0.vernier_delay_line_0.start_pos.n8 tdc_0.vernier_delay_line_0.start_pos.n7 5.74235
R8564 tdc_0.vernier_delay_line_0.start_pos.n13 tdc_0.vernier_delay_line_0.start_pos.n12 5.49235
R8565 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_pos.n13 1.32081
R8566 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_pos.n8 0.40675
R8567 ui_in[7].n0 ui_in[7].t5 628.097
R8568 ui_in[7].n1 ui_in[7].t7 622.766
R8569 ui_in[7].n5 ui_in[7].t2 543.053
R8570 ui_in[7].n0 ui_in[7].t1 523.774
R8571 ui_in[7].n2 ui_in[7].t4 304.647
R8572 ui_in[7].n2 ui_in[7].t6 304.647
R8573 ui_in[7].n5 ui_in[7].t3 221.72
R8574 ui_in[7].n6 ui_in[7].n5 220.327
R8575 ui_in[7].n2 ui_in[7].t0 202.44
R8576 ui_in[7] ui_in[7].n2 169.071
R8577 ui_in[7] ui_in[7].n1 166.244
R8578 ui_in[7].n4 ui_in[7] 35.9653
R8579 ui_in[7].n4 ui_in[7].n3 3.04693
R8580 ui_in[7].n3 ui_in[7] 1.24128
R8581 ui_in[7].n1 ui_in[7].n0 1.09595
R8582 ui_in[7].n3 ui_in[7] 0.402286
R8583 ui_in[7].n6 ui_in[7] 0.063
R8584 ui_in[7] ui_in[7].n4 0.0505
R8585 ui_in[7] ui_in[7].n6 0.0433571
R8586 ui_in[6].n0 ui_in[6].t1 628.097
R8587 ui_in[6].n1 ui_in[6].t5 622.766
R8588 ui_in[6].n5 ui_in[6].t2 543.053
R8589 ui_in[6].n0 ui_in[6].t0 523.774
R8590 ui_in[6].n2 ui_in[6].t7 304.647
R8591 ui_in[6].n2 ui_in[6].t4 304.647
R8592 ui_in[6].n5 ui_in[6].t3 221.72
R8593 ui_in[6].n6 ui_in[6].n5 220.327
R8594 ui_in[6].n2 ui_in[6].t6 202.44
R8595 ui_in[6] ui_in[6].n2 169.071
R8596 ui_in[6] ui_in[6].n1 166.244
R8597 ui_in[6].n4 ui_in[6] 33.1777
R8598 ui_in[6].n4 ui_in[6].n3 2.26836
R8599 ui_in[6].n3 ui_in[6] 1.24128
R8600 ui_in[6].n1 ui_in[6].n0 1.09595
R8601 ui_in[6] ui_in[6].n4 0.761214
R8602 ui_in[6].n3 ui_in[6] 0.402286
R8603 ui_in[6] ui_in[6].n6 0.111214
R8604 ui_in[6].n6 ui_in[6] 0.063
R8605 uio_in[6].n1 uio_in[6].t3 618.668
R8606 uio_in[6].n0 uio_in[6].t2 618.668
R8607 uio_in[6].n1 uio_in[6].t1 456.997
R8608 uio_in[6].n0 uio_in[6].t0 456.997
R8609 uio_in[6] uio_in[6].n1 161.375
R8610 uio_in[6] uio_in[6].n0 161.375
R8611 uio_in[6].n2 uio_in[6] 38.2853
R8612 uio_in[6] uio_in[6].n2 20.1497
R8613 uio_in[6].n2 uio_in[6] 13.5655
R8614 uio_in[0].n0 uio_in[0].t5 628.097
R8615 uio_in[0].n1 uio_in[0].t7 622.766
R8616 uio_in[0].n5 uio_in[0].t3 543.053
R8617 uio_in[0].n0 uio_in[0].t1 523.774
R8618 uio_in[0].n2 uio_in[0].t2 304.647
R8619 uio_in[0].n2 uio_in[0].t6 304.647
R8620 uio_in[0].n5 uio_in[0].t4 221.72
R8621 uio_in[0].n6 uio_in[0].n5 220.327
R8622 uio_in[0].n2 uio_in[0].t0 202.44
R8623 uio_in[0] uio_in[0].n2 169.071
R8624 uio_in[0] uio_in[0].n1 166.244
R8625 uio_in[0].n4 uio_in[0] 38.2949
R8626 uio_in[0].n4 uio_in[0].n3 3.06836
R8627 uio_in[0].n3 uio_in[0] 1.24128
R8628 uio_in[0].n1 uio_in[0].n0 1.09595
R8629 uio_in[0].n3 uio_in[0] 0.402286
R8630 uio_in[0].n6 uio_in[0] 0.063
R8631 uio_in[0] uio_in[0].n4 0.0469286
R8632 uio_in[0] uio_in[0].n6 0.0255
R8633 tdc_0.vernier_delay_line_0.start_neg.n2 tdc_0.vernier_delay_line_0.start_neg.t14 539.841
R8634 tdc_0.vernier_delay_line_0.start_neg.n1 tdc_0.vernier_delay_line_0.start_neg.t8 539.841
R8635 tdc_0.vernier_delay_line_0.start_neg.n5 tdc_0.vernier_delay_line_0.start_neg.t11 539.841
R8636 tdc_0.vernier_delay_line_0.start_neg.n4 tdc_0.vernier_delay_line_0.start_neg.t12 539.841
R8637 tdc_0.vernier_delay_line_0.start_neg.n2 tdc_0.vernier_delay_line_0.start_neg.t13 215.293
R8638 tdc_0.vernier_delay_line_0.start_neg.n1 tdc_0.vernier_delay_line_0.start_neg.t15 215.293
R8639 tdc_0.vernier_delay_line_0.start_neg.n5 tdc_0.vernier_delay_line_0.start_neg.t9 215.293
R8640 tdc_0.vernier_delay_line_0.start_neg.n4 tdc_0.vernier_delay_line_0.start_neg.t10 215.293
R8641 tdc_0.vernier_delay_line_0.start_neg.n7 tdc_0.vernier_delay_line_0.start_neg.n3 166.144
R8642 tdc_0.vernier_delay_line_0.start_neg.n7 tdc_0.vernier_delay_line_0.start_neg.n6 165.8
R8643 tdc_0.vernier_delay_line_0.start_neg.n0 tdc_0.vernier_delay_line_0.start_neg.t1 85.2499
R8644 tdc_0.vernier_delay_line_0.start_neg.n11 tdc_0.vernier_delay_line_0.start_neg.t7 85.2499
R8645 tdc_0.vernier_delay_line_0.start_neg.n11 tdc_0.vernier_delay_line_0.start_neg.t2 83.7172
R8646 tdc_0.vernier_delay_line_0.start_neg.n0 tdc_0.vernier_delay_line_0.start_neg.t0 83.7172
R8647 tdc_0.vernier_delay_line_0.start_neg.n10 tdc_0.vernier_delay_line_0.start_neg.n8 75.7282
R8648 tdc_0.vernier_delay_line_0.start_neg.n10 tdc_0.vernier_delay_line_0.start_neg.n9 66.3172
R8649 tdc_0.vernier_delay_line_0.start_neg.n3 tdc_0.vernier_delay_line_0.start_neg.n1 36.1505
R8650 tdc_0.vernier_delay_line_0.start_neg.n6 tdc_0.vernier_delay_line_0.start_neg.n4 36.1505
R8651 tdc_0.vernier_delay_line_0.start_neg.n3 tdc_0.vernier_delay_line_0.start_neg.n2 34.5438
R8652 tdc_0.vernier_delay_line_0.start_neg.n6 tdc_0.vernier_delay_line_0.start_neg.n5 34.5438
R8653 tdc_0.vernier_delay_line_0.start_neg.n9 tdc_0.vernier_delay_line_0.start_neg.t3 17.4005
R8654 tdc_0.vernier_delay_line_0.start_neg.n9 tdc_0.vernier_delay_line_0.start_neg.t4 17.4005
R8655 tdc_0.vernier_delay_line_0.start_neg.n8 tdc_0.vernier_delay_line_0.start_neg.t5 9.52217
R8656 tdc_0.vernier_delay_line_0.start_neg.n8 tdc_0.vernier_delay_line_0.start_neg.t6 9.52217
R8657 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n0 6.45821
R8658 tdc_0.vernier_delay_line_0.start_neg.n12 tdc_0.vernier_delay_line_0.start_neg.n10 5.30824
R8659 tdc_0.vernier_delay_line_0.start_neg.n12 tdc_0.vernier_delay_line_0.start_neg.n11 4.94887
R8660 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n7 0.754406
R8661 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n12 0.160656
R8662 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 784.053
R8663 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 784.053
R8664 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 784.053
R8665 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 784.053
R8666 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 539.841
R8667 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 539.841
R8668 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 539.841
R8669 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 539.841
R8670 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 215.293
R8671 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 215.293
R8672 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 215.293
R8673 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 215.293
R8674 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 168.659
R8675 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 167.992
R8676 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 166.144
R8677 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 165.8
R8678 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 85.2499
R8679 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 85.2499
R8680 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 83.7172
R8681 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 83.7172
R8682 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 75.7282
R8683 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 66.3172
R8684 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 36.1505
R8685 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 36.1505
R8686 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 34.5438
R8687 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 34.5438
R8688 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 17.4005
R8689 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 17.4005
R8690 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 17.2391
R8691 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 9.52217
R8692 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 9.52217
R8693 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 6.39571
R8694 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 5.30824
R8695 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 4.94887
R8696 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 1.48097
R8697 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 1.06691
R8698 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.539562
R8699 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.391125
R8700 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 0.160656
R8701 a_10108_33108.n2 a_10108_33108.n1 34.9195
R8702 a_10108_33108.n2 a_10108_33108.n0 25.5407
R8703 a_10108_33108.n3 a_10108_33108.n2 25.2907
R8704 a_10108_33108.n1 a_10108_33108.t3 5.8005
R8705 a_10108_33108.n1 a_10108_33108.t5 5.8005
R8706 a_10108_33108.n0 a_10108_33108.t1 5.8005
R8707 a_10108_33108.n0 a_10108_33108.t0 5.8005
R8708 a_10108_33108.n3 a_10108_33108.t2 5.8005
R8709 a_10108_33108.t4 a_10108_33108.n3 5.8005
R8710 variable_delay_dummy_0.variable_delay_unit_1.in.n0 variable_delay_dummy_0.variable_delay_unit_1.in.t4 607.409
R8711 variable_delay_dummy_0.variable_delay_unit_1.in.n2 variable_delay_dummy_0.variable_delay_unit_1.in.t3 543.053
R8712 variable_delay_dummy_0.variable_delay_unit_1.in.n0 variable_delay_dummy_0.variable_delay_unit_1.in.t5 321.423
R8713 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n2 221.778
R8714 variable_delay_dummy_0.variable_delay_unit_1.in.n2 variable_delay_dummy_0.variable_delay_unit_1.in.t2 221.72
R8715 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n0 161.72
R8716 variable_delay_dummy_0.variable_delay_unit_1.in.n1 variable_delay_dummy_0.variable_delay_unit_1.in.t1 84.7227
R8717 variable_delay_dummy_0.variable_delay_unit_1.in.n1 variable_delay_dummy_0.variable_delay_unit_1.in.t0 84.0867
R8718 variable_delay_dummy_0.variable_delay_unit_1.in.n3 variable_delay_dummy_0.variable_delay_unit_1.in 20.0791
R8719 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n3 0.851271
R8720 variable_delay_dummy_0.variable_delay_unit_1.in.n3 variable_delay_dummy_0.variable_delay_unit_1.in.n1 0.465495
R8721 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 variable_delay_dummy_0.variable_delay_unit_1.forward.t2 607.409
R8722 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 variable_delay_dummy_0.variable_delay_unit_1.forward.t3 321.423
R8723 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.forward.n0 161.72
R8724 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 84.7227
R8725 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 84.0867
R8726 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 variable_delay_dummy_0.variable_delay_unit_1.forward 19.7898
R8727 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.forward.n2 0.851271
R8728 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 0.465495
R8729 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 85.1574
R8730 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 83.8097
R8731 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 74.288
R8732 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 67.7574
R8733 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 17.4005
R8734 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 17.4005
R8735 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 9.52217
R8736 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 9.52217
R8737 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 5.83219
R8738 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 5.49235
R8739 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 1.32081
R8740 ui_in[2].n0 ui_in[2].t0 577.653
R8741 ui_in[2].n0 ui_in[2] 37.1928
R8742 ui_in[2] ui_in[2].n0 0.0747188
R8743 uo_out[1].n0 uo_out[1].t4 734.539
R8744 uo_out[1].n0 uo_out[1].t5 233.26
R8745 uo_out[1].n2 uo_out[1].n0 162.335
R8746 uo_out[1].n2 uo_out[1].n1 75.5733
R8747 uo_out[1].n4 uo_out[1].n3 66.3172
R8748 uo_out[1].n5 uo_out[1] 30.7309
R8749 uo_out[1].n3 uo_out[1].t2 17.4005
R8750 uo_out[1].n3 uo_out[1].t0 17.4005
R8751 uo_out[1].n1 uo_out[1].t1 9.52217
R8752 uo_out[1].n1 uo_out[1].t3 9.52217
R8753 uo_out[1].n5 uo_out[1].n4 5.02496
R8754 uo_out[1].n4 uo_out[1].n2 0.438
R8755 uo_out[1] uo_out[1].n5 0.063
R8756 uo_out[2].n0 uo_out[2].t4 734.539
R8757 uo_out[2].n0 uo_out[2].t5 233.26
R8758 uo_out[2].n2 uo_out[2].n0 162.335
R8759 uo_out[2].n2 uo_out[2].n1 75.5733
R8760 uo_out[2].n4 uo_out[2].n3 66.3172
R8761 uo_out[2].n5 uo_out[2] 27.8652
R8762 uo_out[2].n3 uo_out[2].t0 17.4005
R8763 uo_out[2].n3 uo_out[2].t2 17.4005
R8764 uo_out[2].n1 uo_out[2].t3 9.52217
R8765 uo_out[2].n1 uo_out[2].t1 9.52217
R8766 uo_out[2].n5 uo_out[2].n4 5.02496
R8767 uo_out[2].n4 uo_out[2].n2 0.438
R8768 uo_out[2] uo_out[2].n5 0.063
R8769 uio_in[3].n0 uio_in[3].t0 577.653
R8770 uio_in[3].n0 uio_in[3] 39.6907
R8771 uio_in[3] uio_in[3].n0 0.0747188
R8772 ui_in[0].n0 ui_in[0].t0 577.653
R8773 ui_in[0].n0 ui_in[0] 40.4285
R8774 ui_in[0] ui_in[0].n0 0.0747188
R8775 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 890.727
R8776 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 742.783
R8777 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 641.061
R8778 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 623.388
R8779 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 547.874
R8780 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 431.807
R8781 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 427.875
R8782 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 340.632
R8783 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 208.631
R8784 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 168.007
R8785 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R8786 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R8787 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R8788 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R8789 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R8790 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 8.91506
R8791 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R8792 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R8793 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R8794 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R8795 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 879.481
R8796 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 742.783
R8797 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 641.061
R8798 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 623.388
R8799 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 547.874
R8800 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 431.807
R8801 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 427.875
R8802 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 333.161
R8803 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 208.668
R8804 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 168.077
R8805 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R8806 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R8807 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R8808 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 11.1806
R8809 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 10.4291
R8810 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8811 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R8812 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 0.740618
R8813 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 0.228761
R8814 a_10108_37672.n3 a_10108_37672.n2 34.9195
R8815 a_10108_37672.n2 a_10108_37672.n1 25.5407
R8816 a_10108_37672.n2 a_10108_37672.n0 25.2907
R8817 a_10108_37672.n1 a_10108_37672.t0 5.8005
R8818 a_10108_37672.n1 a_10108_37672.t1 5.8005
R8819 a_10108_37672.n0 a_10108_37672.t2 5.8005
R8820 a_10108_37672.n0 a_10108_37672.t5 5.8005
R8821 a_10108_37672.n3 a_10108_37672.t3 5.8005
R8822 a_10108_37672.t4 a_10108_37672.n3 5.8005
R8823 ua[0].n14 ua[0].n13 1348.04
R8824 ua[0].n3 ua[0].n2 1307.92
R8825 ua[0].n5 ua[0].n2 551.179
R8826 ua[0].n16 ua[0].n13 485.663
R8827 ua[0].n19 ua[0].n11 143.792
R8828 ua[0].n19 ua[0].n18 143.792
R8829 ua[0].n7 ua[0].n0 139.512
R8830 ua[0].n7 ua[0].n6 139.512
R8831 ua[0].n1 ua[0].t3 84.7934
R8832 ua[0].n21 ua[0].t4 84.7879
R8833 ua[0].n12 ua[0].t1 84.7879
R8834 ua[0].n4 ua[0].t2 57.2869
R8835 ua[0].n7 ua[0].n2 46.2505
R8836 ua[0].n15 ua[0].t0 44.5923
R8837 ua[0].n18 ua[0].n16 33.509
R8838 ua[0].n6 ua[0].n5 32.2656
R8839 ua[0].n3 ua[0].n0 20.5561
R8840 ua[0].n4 ua[0].n3 20.5561
R8841 ua[0].n14 ua[0].n11 20.5561
R8842 ua[0].n15 ua[0].n14 20.5561
R8843 ua[0].n19 ua[0].n13 18.5005
R8844 ua[0].n17 ua[0] 14.3934
R8845 ua[0].n5 ua[0].n4 8.66346
R8846 ua[0].n16 ua[0].n15 7.4066
R8847 ua[0].n8 ua[0].n7 2.3255
R8848 ua[0].n9 ua[0].n0 2.2281
R8849 ua[0].n6 ua[0].n1 2.17472
R8850 ua[0].n22 ua[0].n11 2.0406
R8851 ua[0].n18 ua[0].n17 2.0406
R8852 ua[0].n20 ua[0].n19 1.8605
R8853 ua[0] ua[0].n10 0.620598
R8854 ua[0].n10 ua[0].n9 0.223
R8855 ua[0].n22 ua[0].n21 0.129176
R8856 ua[0].n17 ua[0].n12 0.124275
R8857 ua[0].n20 ua[0].n12 0.110794
R8858 ua[0].n21 ua[0].n20 0.105892
R8859 ua[0].n8 ua[0].n1 0.0577917
R8860 ua[0] ua[0].n22 0.0103039
R8861 ua[0].n10 ua[0] 0.00540196
R8862 ua[0].n9 ua[0].n8 0.00440625
R8863 variable_delay_short_0.variable_delay_unit_2.in.n0 variable_delay_short_0.variable_delay_unit_2.in.t5 607.409
R8864 variable_delay_short_0.variable_delay_unit_2.in.n2 variable_delay_short_0.variable_delay_unit_2.in.t2 543.053
R8865 variable_delay_short_0.variable_delay_unit_2.in.n0 variable_delay_short_0.variable_delay_unit_2.in.t4 321.423
R8866 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n2 221.778
R8867 variable_delay_short_0.variable_delay_unit_2.in.n2 variable_delay_short_0.variable_delay_unit_2.in.t3 221.72
R8868 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n0 161.72
R8869 variable_delay_short_0.variable_delay_unit_2.in.n1 variable_delay_short_0.variable_delay_unit_2.in.t0 84.7227
R8870 variable_delay_short_0.variable_delay_unit_2.in.n1 variable_delay_short_0.variable_delay_unit_2.in.t1 84.0867
R8871 variable_delay_short_0.variable_delay_unit_2.in.n3 variable_delay_short_0.variable_delay_unit_2.in 20.0791
R8872 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n3 0.851271
R8873 variable_delay_short_0.variable_delay_unit_2.in.n3 variable_delay_short_0.variable_delay_unit_2.in.n1 0.465495
R8874 variable_delay_short_0.variable_delay_unit_1.in.n0 variable_delay_short_0.variable_delay_unit_1.in.t5 607.409
R8875 variable_delay_short_0.variable_delay_unit_1.in.n2 variable_delay_short_0.variable_delay_unit_1.in.t2 543.053
R8876 variable_delay_short_0.variable_delay_unit_1.in.n0 variable_delay_short_0.variable_delay_unit_1.in.t4 321.423
R8877 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n2 221.778
R8878 variable_delay_short_0.variable_delay_unit_1.in.n2 variable_delay_short_0.variable_delay_unit_1.in.t3 221.72
R8879 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n0 161.72
R8880 variable_delay_short_0.variable_delay_unit_1.in.n1 variable_delay_short_0.variable_delay_unit_1.in.t1 84.7227
R8881 variable_delay_short_0.variable_delay_unit_1.in.n1 variable_delay_short_0.variable_delay_unit_1.in.t0 84.0867
R8882 variable_delay_short_0.variable_delay_unit_1.in.n3 variable_delay_short_0.variable_delay_unit_1.in 20.0791
R8883 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n3 0.851271
R8884 variable_delay_short_0.variable_delay_unit_1.in.n3 variable_delay_short_0.variable_delay_unit_1.in.n1 0.465495
R8885 ui_in[3].n0 ui_in[3].t0 727.072
R8886 ui_in[3].n0 ui_in[3] 36.9161
R8887 ui_in[3].n0 ui_in[3] 0.323417
R8888 ui_in[3] ui_in[3].n0 0.0610469
R8889 uio_in[1].n0 uio_in[1].t0 577.653
R8890 uio_in[1].n0 uio_in[1] 42.0234
R8891 uio_in[1] uio_in[1].n0 0.0747188
R8892 uio_in[4].n0 uio_in[4].t0 727.072
R8893 uio_in[4].n0 uio_in[4] 39.7322
R8894 uio_in[4].n0 uio_in[4] 0.323417
R8895 uio_in[4] uio_in[4].n0 0.0610469
R8896 uio_in[5].n0 uio_in[5].t1 564.04
R8897 uio_in[5].n0 uio_in[5].t0 511.623
R8898 uio_in[5].n1 uio_in[5].n0 161.3
R8899 uio_in[5].n1 uio_in[5] 50.8219
R8900 uio_in[5] uio_in[5].n1 0.0295179
R8901 ui_in[1].n0 ui_in[1].t0 727.072
R8902 ui_in[1].n0 ui_in[1] 40.1518
R8903 ui_in[1].n0 ui_in[1] 0.323417
R8904 ui_in[1] ui_in[1].n0 0.0610469
R8905 uio_in[2].n0 uio_in[2].t0 727.072
R8906 uio_in[2].n0 uio_in[2] 42.3292
R8907 uio_in[2].n0 uio_in[2] 0.323417
R8908 uio_in[2] uio_in[2].n0 0.0610469
C0 input_stage_andpwr_0.fine_delay_unit_1.in ui_in[1] 0.039118f
C1 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[6] 9.38e-20
C2 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.forward 7.91e-21
C3 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.in 8.82e-20
C4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 8.54e-19
C5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.start_pos 4.53e-19
C6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_13254_37444# 0.010872f
C7 a_12310_30552# a_13254_30598# 1.02e-19
C8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_13254_28316# 0.010872f
C9 input_stage_andpwr_0.fine_delay_unit_0.in a_24790_6672# 0.244525f
C10 variable_delay_short_0.out uio_in[3] 0.036391f
C11 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 6.08e-20
C12 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.in 0.09141f
C13 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.192064f
C14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 uo_out[2] 3.69e-19
C15 a_12310_32834# uo_out[4] 0.098308f
C16 a_24240_14314# ui_in[7] 0.042718f
C17 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C18 variable_delay_short_0.variable_delay_unit_4.out a_25060_21092# 0.070146f
C19 a_12420_33258# VDPWR 0.497547f
C20 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.in 8.82e-20
C21 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12308_28732# 3.26e-19
C22 VDPWR a_15680_11634# 1.70112f
C23 variable_delay_short_0.variable_delay_unit_2.out ui_in[5] 2.67e-19
C24 input_stage_0.fine_delay_unit_1.in uio_in[6] 1.82e-20
C25 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12420_39726# 0.003664f
C26 VDPWR a_13254_28316# 6.18e-19
C27 a_9330_15214# a_9330_15794# 0.001101f
C28 a_25060_23158# ui_in[2] 3.98e-20
C29 a_12420_26034# a_12310_25988# 0.030392f
C30 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.out 0.172055f
C31 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VDPWR 2.55561f
C32 a_12420_33258# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.033952f
C33 a_15680_11634# variable_delay_dummy_0.in 8.82e-20
C34 variable_delay_short_0.variable_delay_unit_1.in ui_in[3] 0.02f
C35 VDPWR uo_out[7] 0.587468f
C36 uio_in[3] uio_in[1] 0.001793f
C37 a_10108_25734# a_12310_25988# 2.08e-21
C38 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_12420_28316# 1.47e-19
C39 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.010157f
C40 variable_delay_short_0.variable_delay_unit_3.in ui_in[7] 3.37e-20
C41 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.231672f
C42 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VDPWR 0.706489f
C43 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 1.24e-19
C44 uio_oe[3] uio_oe[2] 0.170937f
C45 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.100263f
C46 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[2] 6.97e-19
C47 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[2] 2.77e-19
C48 a_12310_37398# uo_out[6] 0.098308f
C49 a_12308_31014# uo_out[4] 6.49e-20
C50 a_24790_6672# input_stage_andpwr_0.nand_gate_0.out 5.26e-20
C51 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.100263f
C52 input_stage_0.fine_delay_unit_0.in uio_in[6] 6.7e-20
C53 ui_in[7] ui_in[3] 0.014973f
C54 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 1.24e-19
C55 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.53e-19
C56 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.vernier_delay_line_0.start_neg 0.036472f
C57 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en ui_in[6] 1.09842f
C58 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.2373f
C59 a_25060_20210# ui_in[5] 0.15982f
C60 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 uo_out[1] 1.53e-22
C61 VDPWR uo_out[1] 0.587468f
C62 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 5.07283f
C63 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12310_23706# 0.014814f
C64 variable_delay_short_0.variable_delay_unit_4.out VDPWR 1.3445f
C65 a_24240_24040# ui_in[5] 2.89e-20
C66 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.752988f
C67 variable_delay_short_0.variable_delay_unit_4.in a_24240_21092# 0.020173f
C68 a_25060_26988# ui_in[4] 8.92e-19
C69 a_9330_15214# tdc_0.diff_gen_0.delay_unit_2_2.in_2 5.93e-19
C70 a_12420_35540# uo_out[5] 0.013457f
C71 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 a_10108_34862# 0.007929f
C72 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 1.06381f
C73 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 6.93e-19
C74 a_12420_35540# a_13254_35540# 0.003413f
C75 VDPWR ui_in[6] 1.41131f
C76 variable_delay_short_0.variable_delay_unit_3.out ui_in[5] 0.22469f
C77 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_10108_39426# 1.06381f
C78 a_25060_21092# ui_in[2] 3.98e-20
C79 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_16500_12516# 0.15982f
C80 variable_delay_dummy_0.variable_delay_unit_1.out VDPWR 1.61031f
C81 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.forward 0.016896f
C82 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_24240_24040# 0.029284f
C83 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12420_23752# 0.035356f
C84 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 1.24e-19
C85 input_stage_andpwr_0.nand_gate_0.out a_25284_5108# 0.355469f
C86 a_12310_28270# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 6.08e-20
C87 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_12310_32834# 3.84e-19
C88 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.007929f
C89 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[6] 0.10528f
C90 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[2] 6.28e-22
C91 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 uo_out[1] 0.20241f
C92 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.45e-19
C93 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.out 0.12029f
C94 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 8.54e-19
C95 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en ui_in[4] 9.38e-20
C96 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.vernier_delay_line_0.start_neg 0.286409f
C97 a_24240_15196# a_25060_15196# 0.011184f
C98 a_12308_35578# a_12310_35116# 0.00595f
C99 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35162# 0.013457f
C100 a_25060_26106# ui_in[3] 0.002391f
C101 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.out 0.002141f
C102 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.in 0.087283f
C103 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 uo_out[3] 1.53e-22
C104 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en ui_in[2] 6.97e-19
C105 a_24790_8314# ui_in[2] 0.024917f
C106 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C107 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.311186f
C108 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_delay 1.12095f
C109 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 8.54e-19
C110 uo_out[7] uo_out[6] 0.856749f
C111 a_25060_23158# VDPWR 6.98e-19
C112 a_9330_14054# variable_delay_short_0.out 7.21e-19
C113 a_15680_14582# uio_in[6] 0.001509f
C114 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_15680_15464# 0.029284f
C115 a_12308_26450# uo_out[1] 0.014835f
C116 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq uo_out[2] 0.229249f
C117 a_12420_32880# VDPWR 0.497771f
C118 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.57093f
C119 tdc_0.diff_gen_0.delay_unit_2_1.in_2 VDPWR 3.06163f
C120 VDPWR a_24240_11366# 1.6584f
C121 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 1.17e-19
C122 VDPWR ui_in[2] 0.001157f
C123 a_13254_24130# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.012202f
C124 a_13254_24130# VDPWR 6.18e-19
C125 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 5.20504f
C126 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.138497f
C127 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.953579f
C128 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37822# 0.504416f
C129 a_12308_37860# a_13254_37822# 1.02e-19
C130 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[4] 0.025512f
C131 a_12310_25988# a_13254_26034# 1.02e-19
C132 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.006183f
C133 uo_out[5] uo_out[2] 2.26e-21
C134 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en VDPWR 2.77611f
C135 uo_out[4] uo_out[3] 1.91867f
C136 a_12308_28732# a_13254_28694# 1.02e-19
C137 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28694# 0.504416f
C138 a_12420_32880# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.003664f
C139 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.747722f
C140 a_12420_32880# a_13254_32880# 0.003413f
C141 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 6.79e-20
C142 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out 0.071795f
C143 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq uo_out[0] 0.229249f
C144 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12308_35578# 0.197073f
C145 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 uo_out[1] 0.10528f
C146 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[4] 4.58e-20
C147 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 3.23832f
C148 input_stage_andpwr_0.fine_delay_unit_1.in ui_in[2] 0.010002f
C149 a_12310_23706# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 3.84e-19
C150 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.871529f
C151 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.283838f
C152 uo_out[1] uo_out[0] 2.98059f
C153 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.018644f
C154 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.756572f
C155 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_12310_25988# 3.84e-19
C156 a_13254_40104# uo_out[7] 0.005712f
C157 variable_delay_short_0.variable_delay_unit_1.out uio_in[0] 0.043504f
C158 a_25060_21092# VDPWR 0.001468f
C159 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 4.53e-19
C160 variable_delay_dummy_0.variable_delay_unit_1.forward a_15680_14582# 0.088132f
C161 variable_delay_short_0.variable_delay_unit_4.out ui_in[5] 0.043597f
C162 a_9330_15214# a_9330_14924# 0.083149f
C163 variable_delay_dummy_0.variable_delay_unit_1.out a_15680_12516# 0.071074f
C164 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12310_30552# 0.196592f
C165 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 uo_out[5] 1.35e-20
C166 a_12310_32834# a_12308_31014# 0.005984f
C167 a_12420_35162# uo_out[5] 0.492009f
C168 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_24240_20210# 0.11539f
C169 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 1.24e-19
C170 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.752988f
C171 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.132512f
C172 a_24240_24040# variable_delay_short_0.variable_delay_unit_5.in 0.020173f
C173 a_15680_11634# uio_in[5] 0.002316f
C174 a_25060_26988# ui_in[3] 0.002391f
C175 ua[0] ui_in[1] 0.002217f
C176 ui_in[5] ui_in[6] 5.05846f
C177 a_16500_11634# uio_in[2] 3.05e-20
C178 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.132512f
C179 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward 0.234428f
C180 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.out 0.12029f
C181 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_13254_23752# 0.010872f
C182 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 a_12310_37398# 3.84e-19
C183 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq uo_out[7] 0.229856f
C184 VDPWR variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 2.77611f
C185 a_9330_14344# variable_delay_short_0.out 3.54e-19
C186 variable_delay_short_0.out a_25060_12248# 0.172055f
C187 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.57093f
C188 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 1.24e-19
C189 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[3] 0.00127f
C190 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.in 0.09141f
C191 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en ui_in[6] 2.92e-19
C192 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.out 0.172055f
C193 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35162# 0.005542f
C194 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_25060_11366# 2.39e-19
C195 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en ui_in[3] 0.014554f
C196 a_24790_6936# ui_in[1] 0.024305f
C197 a_13254_28694# uo_out[2] 0.005542f
C198 a_12420_26412# uo_out[1] 0.013457f
C199 a_23820_8460# a_24790_8050# 0.53267f
C200 input_stage_andpwr_0.fine_delay_unit_1.in a_24790_8314# 0.028846f
C201 a_24240_18144# a_25060_18144# 0.011184f
C202 a_25060_11366# variable_delay_short_0.in 8.82e-20
C203 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 2.43941f
C204 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 3.23844f
C205 a_12420_37822# a_13254_37822# 0.003413f
C206 a_24240_15196# ui_in[3] 0.001719f
C207 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.93e-19
C208 variable_delay_dummy_0.out a_15680_11634# 0.505512f
C209 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.441213f
C210 a_9330_14924# tdc_0.diff_gen_0.delay_unit_2_1.in_1 2.18e-19
C211 a_23820_8460# variable_delay_short_0.in 0.121301f
C212 a_25060_12248# uio_in[0] 0.001909f
C213 a_12420_28694# a_13254_28694# 0.003413f
C214 a_12310_37398# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 6.08e-20
C215 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.28924f
C216 a_13254_24130# uo_out[0] 0.005542f
C217 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12420_35540# 0.033952f
C218 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.out 0.12029f
C219 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 uo_out[0] 1.35e-20
C220 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 2.43248f
C221 variable_delay_short_0.variable_delay_unit_5.forward ui_in[4] 0.036352f
C222 a_13254_32880# VDPWR 6.18e-19
C223 VDPWR variable_delay_dummy_0.in 1.61964f
C224 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 3.6e-19
C225 a_12310_23706# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.164402f
C226 ui_in[5] ui_in[2] 7.13e-19
C227 a_12310_23706# VDPWR 1.42748f
C228 input_stage_andpwr_0.fine_delay_unit_1.in VDPWR 1.33496f
C229 VDPWR tdc_0.diff_gen_0.delay_unit_2_3.in_2 3.06075f
C230 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.138497f
C231 a_12310_23706# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 4.55e-19
C232 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.019931f
C233 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37444# 0.013457f
C234 a_12308_37860# a_12310_37398# 0.00595f
C235 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 2.59e-20
C236 a_25284_5108# uio_in[6] 0.009499f
C237 a_12308_28732# a_12310_28270# 0.00595f
C238 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28316# 0.013457f
C239 input_stage_andpwr_0.fine_delay_unit_0.in ui_in[1] 0.021403f
C240 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_12310_25988# 4.55e-19
C241 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.15e-21
C242 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_25060_23158# 2.39e-19
C243 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 uo_out[4] 0.20241f
C244 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.871529f
C245 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[3] 0.014554f
C246 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[5] 0.016377f
C247 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 2.57093f
C248 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 4.53e-19
C249 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 6.79e-20
C250 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.006183f
C251 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.59e-20
C252 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en ui_in[2] 6.97e-19
C253 variable_delay_dummy_0.variable_delay_unit_1.in uio_in[2] 1.1e-20
C254 a_9330_15504# VDPWR 1.1544f
C255 a_12420_23752# a_13254_23752# 0.003413f
C256 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VDPWR 1.93357f
C257 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12310_39680# 0.196592f
C258 variable_delay_short_0.variable_delay_unit_1.out a_24240_12248# 0.071074f
C259 a_25060_15196# variable_delay_short_0.variable_delay_unit_2.out 0.070146f
C260 variable_delay_short_0.out ui_in[1] 0.001119f
C261 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 uo_out[5] 3.69e-19
C262 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12308_26450# 7.19e-22
C263 a_12308_33296# uo_out[5] 6.49e-20
C264 a_12310_39680# uo_out[7] 0.098487f
C265 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.283838f
C266 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.871529f
C267 variable_delay_short_0.variable_delay_unit_3.in a_24240_18144# 0.020173f
C268 a_24240_24040# variable_delay_short_0.variable_delay_unit_5.out 0.071074f
C269 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_10108_34862# 1.06381f
C270 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDPWR 0.706518f
C271 VDPWR a_15322_8490# 1.25073f
C272 a_24240_18144# ui_in[3] 0.001719f
C273 a_25060_21092# ui_in[5] 0.001909f
C274 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 a_12310_37398# 4.55e-19
C275 tdc_0.start_buffer_0.start_buff a_7140_10670# 0.684455f
C276 VDPWR uio_in[4] 0.004419f
C277 VDPWR tdc_0.diff_gen_0.delay_unit_2_3.in_1 4.44087f
C278 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.in 0.091118f
C279 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out 0.071795f
C280 a_24790_8050# variable_delay_short_0.in 3.44e-20
C281 VDPWR a_12308_26450# 1.40782f
C282 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.79e-20
C283 input_stage_andpwr_0.nand_gate_0.out ui_in[1] 6.37e-19
C284 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12308_37860# 0.197073f
C285 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12308_28732# 0.197073f
C286 variable_delay_short_0.variable_delay_unit_1.out a_24240_14314# 0.505512f
C287 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 a_12310_35116# 3.84e-19
C288 a_13254_35162# uo_out[5] 0.188081f
C289 a_12420_35162# a_12310_35116# 0.030392f
C290 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.in 0.235667f
C291 variable_delay_short_0.variable_delay_unit_5.out ui_in[1] 0.001119f
C292 variable_delay_dummy_0.in a_15322_8490# 0.123564f
C293 variable_delay_dummy_0.in uio_in[4] 0.03818f
C294 variable_delay_short_0.variable_delay_unit_1.in a_25060_11366# 0.054206f
C295 VDPWR uo_out[6] 0.587468f
C296 uio_out[6] uio_out[7] 0.170937f
C297 variable_delay_short_0.variable_delay_unit_2.in uio_in[0] 3.37e-20
C298 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12308_37860# 7.19e-22
C299 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 2.36e-21
C300 a_15322_7112# VDPWR 1.25441f
C301 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.667766f
C302 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en ui_in[5] 9.38e-20
C303 a_12308_24168# a_12310_25988# 0.005984f
C304 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 1.99e-19
C305 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 2.43248f
C306 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.018644f
C307 variable_delay_short_0.variable_delay_unit_5.in ui_in[6] 0.001598f
C308 a_12308_31014# a_12420_30976# 0.030083f
C309 a_12308_31014# uo_out[3] 0.014835f
C310 a_12308_37860# uo_out[7] 6.49e-20
C311 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 3.84e-19
C312 tdc_0.start_buffer_0.start_buff a_9330_13764# 5.99e-19
C313 VDPWR a_15680_12516# 1.78275f
C314 a_9330_14634# a_9330_14344# 0.083149f
C315 a_24240_24040# ui_in[4] 0.127858f
C316 a_9330_14054# a_9330_15794# 5.08e-20
C317 a_24240_12248# a_25060_12248# 0.011184f
C318 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 uo_out[0] 0.10528f
C319 VDPWR uo_out[0] 0.587468f
C320 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 uo_out[0] 3.69e-19
C321 a_12420_26034# uo_out[1] 0.492009f
C322 a_12310_28270# uo_out[2] 0.098308f
C323 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12308_26450# 0.162625f
C324 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.499806f
C325 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.out 0.172055f
C326 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 VDPWR 2.23953f
C327 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.441213f
C328 uio_oe[2] uio_oe[1] 0.170937f
C329 a_15680_12516# variable_delay_dummy_0.in 7.65e-21
C330 VDPWR ui_in[5] 1.43813f
C331 variable_delay_short_0.variable_delay_unit_3.out ui_in[4] 2.67e-19
C332 variable_delay_short_0.variable_delay_unit_1.out ui_in[3] 0.040959f
C333 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.499806f
C334 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.138497f
C335 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.019931f
C336 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 1.17e-19
C337 a_12310_23706# uo_out[0] 0.098308f
C338 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12420_35162# 0.003664f
C339 VDPWR a_24240_26106# 1.70112f
C340 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 5.04e-20
C341 tdc_0.start_buffer_0.start_buff tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.001356f
C342 uio_out[5] uio_out[4] 0.170937f
C343 a_15322_8490# uio_in[4] 0.010812f
C344 a_16500_11634# uio_in[3] 4.35e-20
C345 a_13254_40104# VDPWR 6.18e-19
C346 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.006183f
C347 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VDPWR 5.07283f
C348 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 4.28924f
C349 a_25060_23158# variable_delay_short_0.variable_delay_unit_5.in 0.054206f
C350 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en VDPWR 2.7762f
C351 variable_delay_dummy_0.variable_delay_unit_1.out a_16500_14582# 0.222585f
C352 variable_delay_short_0.variable_delay_unit_5.forward ui_in[3] 0.007775f
C353 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.in 8.82e-20
C354 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37444# 0.005542f
C355 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28316# 0.005542f
C356 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.010157f
C357 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[5] 6.28e-22
C358 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.138497f
C359 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C360 variable_delay_dummy_0.in a_16292_8080# 3.44e-20
C361 variable_delay_short_0.variable_delay_unit_5.in ui_in[2] 3.31e-20
C362 a_15322_7112# a_15322_8490# 0.001571f
C363 a_13254_30976# VDPWR 6.18e-19
C364 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.814958f
C365 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en VDPWR 3.86972f
C366 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 uo_out[2] 0.10528f
C367 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 0.031607f
C368 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.in 0.08442f
C369 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12420_37822# 0.033952f
C370 VDPWR a_12420_26412# 0.497547f
C371 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_12308_26450# 0.197073f
C372 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en ui_in[7] 9.38e-20
C373 a_24240_14314# a_25060_14314# 0.004142f
C374 a_9330_14054# a_9330_13764# 0.083149f
C375 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDPWR 0.706518f
C376 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12420_28694# 0.033952f
C377 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 a_12310_35116# 4.55e-19
C378 uo_out[7] uo_out[5] 1.56e-19
C379 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.196592f
C380 variable_delay_short_0.variable_delay_unit_2.out a_24240_17262# 0.505512f
C381 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.010157f
C382 a_12308_33296# a_12310_35116# 0.005984f
C383 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.out 0.235667f
C384 variable_delay_short_0.variable_delay_unit_3.out a_25060_18144# 0.070146f
C385 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.132512f
C386 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.out 0.071795f
C387 uio_in[7] uo_out[0] 0.073214f
C388 a_25060_12248# ui_in[3] 0.002391f
C389 VDPWR uio_in[5] 0.925517f
C390 variable_delay_short_0.variable_delay_unit_2.out ui_in[3] 0.040959f
C391 ui_in[6] uio_in[0] 9.78e-19
C392 a_12308_40142# a_12420_40104# 0.030083f
C393 a_9330_14344# a_9330_15794# 1.76e-19
C394 a_24240_20210# a_25060_20210# 0.004142f
C395 a_23820_7082# ui_in[0] 0.003341f
C396 a_12420_30976# uo_out[3] 0.013457f
C397 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 4.55e-19
C398 uo_out[4] uo_out[2] 1.56e-19
C399 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.36e-21
C400 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.in 7.65e-21
C401 a_23820_8460# a_23820_7082# 0.001571f
C402 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12308_35578# 7.19e-22
C403 a_15322_8490# a_16292_8080# 0.53267f
C404 a_12310_35116# a_13254_35162# 1.02e-19
C405 ui_in[6] uio_in[1] 3.03e-19
C406 input_stage_0.fine_delay_unit_1.in a_16292_8344# 0.028846f
C407 variable_delay_dummy_0.in uio_in[5] 0.060059f
C408 a_16292_8344# uio_in[2] 4.3e-19
C409 a_16292_8080# uio_in[4] 0.00799f
C410 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_24240_21092# 0.029284f
C411 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 uo_out[0] 6.28e-22
C412 variable_delay_dummy_0.variable_delay_unit_1.in uio_in[3] 3.5e-20
C413 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12420_26412# 0.003607f
C414 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.2373f
C415 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.99e-19
C416 a_25060_20210# variable_delay_short_0.variable_delay_unit_3.in 8.82e-20
C417 a_25060_14314# ui_in[3] 0.002391f
C418 variable_delay_short_0.out a_24240_11366# 0.505512f
C419 variable_delay_short_0.variable_delay_unit_3.out a_24240_20210# 0.505512f
C420 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30976# 0.174293f
C421 a_10108_30298# a_12310_30552# 2.08e-21
C422 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_10108_37144# 1.06381f
C423 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 7.19e-22
C424 variable_delay_short_0.out ui_in[2] 0.003069f
C425 VDPWR variable_delay_dummy_0.out 1.79065f
C426 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_10108_28016# 1.06381f
C427 a_25060_20210# ui_in[3] 0.002391f
C428 variable_delay_short_0.variable_delay_unit_4.out ui_in[4] 0.227555f
C429 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.441213f
C430 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 3.26e-19
C431 a_24240_14314# variable_delay_short_0.variable_delay_unit_2.in 0.088132f
C432 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_neg 0.688629f
C433 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.out 0.002141f
C434 VDPWR a_24240_26988# 1.78268f
C435 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VDPWR 3.23832f
C436 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 4.28924f
C437 a_13254_26034# uo_out[1] 0.188081f
C438 VDPWR ua[0] 0.762707f
C439 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003768f
C440 a_25060_15196# ui_in[6] 6.99e-20
C441 a_24240_24040# ui_in[3] 0.001719f
C442 a_24240_17262# a_25060_17262# 0.004142f
C443 variable_delay_short_0.variable_delay_unit_3.in a_25060_17262# 0.054206f
C444 variable_delay_dummy_0.out variable_delay_dummy_0.in 0.728538f
C445 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_3.in 0.499092f
C446 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 uo_out[7] 0.105414f
C447 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12310_25988# 3.45e-19
C448 a_15680_15464# uio_in[6] 0.006769f
C449 a_12420_37444# a_12310_37398# 0.030392f
C450 ui_in[4] ui_in[6] 0.002613f
C451 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 1.17e-19
C452 a_24240_11366# uio_in[0] 0.042718f
C453 a_16292_6966# input_stage_0.fine_delay_unit_1.in 5.97e-19
C454 a_12420_28316# a_12310_28270# 0.030392f
C455 a_25060_17262# ui_in[3] 0.002391f
C456 uio_in[0] ui_in[2] 7.13e-19
C457 a_12308_26450# a_12420_26412# 0.030083f
C458 a_16292_6966# uio_in[2] 0.024305f
C459 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.441213f
C460 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 VDPWR 5.07283f
C461 variable_delay_short_0.variable_delay_unit_3.out ui_in[3] 0.040959f
C462 variable_delay_short_0.variable_delay_unit_5.out ui_in[2] 0.002549f
C463 input_stage_0.fine_delay_unit_1.in uio_in[2] 0.039331f
C464 VDPWR variable_delay_short_0.variable_delay_unit_5.in 2.63444f
C465 a_15322_8490# uio_in[5] 0.01196f
C466 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en uio_in[0] 1.5e-19
C467 uio_in[4] uio_in[5] 7.75329f
C468 a_9330_15214# tdc_0.diff_gen_0.delay_unit_2_1.in_1 5.9e-19
C469 ui_in[3] ui_in[1] 0.018155f
C470 a_12310_39680# VDPWR 1.42789f
C471 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.45e-19
C472 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.in 8.82e-20
C473 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 uo_out[1] 1.35e-20
C474 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.in 0.087283f
C475 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en ui_in[5] 8.8e-19
C476 uio_oe[7] uio_oe[6] 0.170937f
C477 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_12420_26412# 0.033952f
C478 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.814958f
C479 variable_delay_short_0.variable_delay_unit_2.in ui_in[3] 0.02f
C480 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_10108_30298# 0.09966f
C481 variable_delay_short_0.variable_delay_unit_1.in ui_in[7] 0.506369f
C482 ui_in[7] uio_in[2] 2.48e-19
C483 input_stage_0.fine_delay_unit_0.in a_16292_6966# 0.028846f
C484 a_12310_37398# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.15e-21
C485 a_15322_7112# a_16292_6702# 0.53267f
C486 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.59e-20
C487 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 1.17e-19
C488 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 uo_out[5] 0.20241f
C489 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.100263f
C490 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.283838f
C491 a_12310_30552# VDPWR 1.42789f
C492 input_stage_0.fine_delay_unit_0.in input_stage_0.fine_delay_unit_1.in 0.029975f
C493 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.706518f
C494 a_24790_6672# ui_in[0] 0.022037f
C495 a_15322_7112# uio_in[5] 0.007103f
C496 input_stage_andpwr_0.fine_delay_unit_1.in a_24790_6936# 5.97e-19
C497 input_stage_0.fine_delay_unit_0.in uio_in[2] 0.021403f
C498 a_25060_23158# ui_in[4] 0.15982f
C499 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.start_buffer_0.start_delay 0.04313f
C500 variable_delay_dummy_0.out a_15322_8490# 0.011089f
C501 a_15680_11634# uio_in[6] 0.001509f
C502 a_25060_15196# ui_in[2] 3.98e-20
C503 VDPWR a_12420_26034# 0.497771f
C504 a_16500_14582# VDPWR 0.160518f
C505 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12420_37444# 0.003664f
C506 a_15680_12516# uio_in[5] 0.002316f
C507 variable_delay_dummy_0.out uio_in[4] 0.007407f
C508 a_24790_8314# variable_delay_short_0.out 4.38e-19
C509 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12420_28316# 0.003664f
C510 uo_out[0] uio_in[5] 1.17e-19
C511 input_stage_andpwr_0.fine_delay_unit_0.in VDPWR 0.323759f
C512 ui_in[4] ui_in[2] 7.13e-19
C513 a_25060_18144# ui_in[6] 0.001909f
C514 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_25060_15196# 0.15982f
C515 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.forward 0.016896f
C516 a_12308_37860# VDPWR 1.40782f
C517 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.747722f
C518 a_16786_5138# VDPWR 0.002853f
C519 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.79e-20
C520 tdc_0.diff_gen_0.delay_unit_2_6.in_2 VDPWR 3.06151f
C521 a_10108_39426# a_12310_39680# 2.08e-21
C522 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_13254_40104# 0.174293f
C523 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_15680_11634# 0.11539f
C524 a_12420_30598# uo_out[3] 0.492009f
C525 input_stage_andpwr_0.fine_delay_unit_1.in input_stage_andpwr_0.fine_delay_unit_0.in 0.029975f
C526 VDPWR variable_delay_short_0.out 1.72578f
C527 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.99e-19
C528 a_16292_8080# uio_in[5] 0.002587f
C529 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 9.61e-20
C530 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C531 a_15680_12516# variable_delay_dummy_0.out 0.493816f
C532 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12420_26034# 0.035356f
C533 a_24240_24040# a_25060_24040# 0.011184f
C534 uo_out[1] uio_in[6] 1.2e-19
C535 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 uo_out[6] 1.35e-20
C536 variable_delay_short_0.out variable_delay_dummy_0.in 0.100566f
C537 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.132512f
C538 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12310_30552# 0.014814f
C539 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.752988f
C540 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.132512f
C541 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C542 input_stage_andpwr_0.fine_delay_unit_1.in variable_delay_short_0.out 0.024792f
C543 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.752988f
C544 input_stage_andpwr_0.nand_gate_0.out VDPWR 0.275003f
C545 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_10108_25734# 1.06381f
C546 a_12308_33296# uo_out[4] 0.014835f
C547 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 VDPWR 3.23832f
C548 a_25060_21092# ui_in[4] 6.99e-20
C549 VDPWR uio_in[0] 1.46811f
C550 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14634# 0.00141f
C551 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.006183f
C552 VDPWR variable_delay_short_0.variable_delay_unit_5.out 1.5668f
C553 a_24240_26988# ui_in[5] 2.89e-20
C554 a_25060_18144# ui_in[2] 3.98e-20
C555 variable_delay_short_0.variable_delay_unit_4.out ui_in[3] 0.040959f
C556 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 uo_out[1] 3.69e-19
C557 tdc_0.diff_gen_0.delay_unit_2_6.in_1 VDPWR 4.42926f
C558 VDPWR uio_in[1] 6.39e-19
C559 a_24240_17262# ui_in[6] 0.042718f
C560 variable_delay_dummy_0.out a_16292_8080# 6.96e-19
C561 variable_delay_short_0.variable_delay_unit_3.in ui_in[6] 0.580889f
C562 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[6] 0.005546f
C563 a_12310_37398# a_13254_37444# 1.02e-19
C564 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.706518f
C565 a_12310_28270# a_13254_28316# 1.02e-19
C566 a_16292_6702# uio_in[5] 9.94e-20
C567 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26412# 0.174293f
C568 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.953579f
C569 ui_in[6] ui_in[3] 0.014973f
C570 a_12308_33296# a_13254_33258# 1.02e-19
C571 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_33258# 0.504416f
C572 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C573 a_15680_15464# a_16500_15464# 0.011184f
C574 variable_delay_short_0.variable_delay_unit_5.in ui_in[5] 0.00265f
C575 a_16292_8344# uio_in[3] 0.025624f
C576 VDPWR uo_out[5] 0.587468f
C577 VDPWR a_13254_35540# 6.18e-19
C578 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_10108_28016# 0.192064f
C579 input_stage_0.nand_gate_0.out VDPWR 1.25731f
C580 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.out 0.002141f
C581 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.085059f
C582 variable_delay_short_0.out a_15322_8490# 7.6e-19
C583 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.in 8.82e-20
C584 tdc_0.start_buffer_0.start_delay VDPWR 4.05162f
C585 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_12420_26034# 0.003664f
C586 a_25060_15196# VDPWR 0.001468f
C587 variable_delay_short_0.out uio_in[4] 0.10432f
C588 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.231672f
C589 a_12308_37860# uo_out[6] 0.014835f
C590 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[5] 1.53e-22
C591 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_24240_14314# 0.11539f
C592 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.in 0.814958f
C593 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12310_35116# 0.196592f
C594 VDPWR ui_in[4] 1.64573f
C595 a_12420_37822# VDPWR 0.497547f
C596 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_10108_25734# 0.09966f
C597 a_12308_28732# uo_out[3] 6.49e-20
C598 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 2.59e-20
C599 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.100263f
C600 VDPWR a_13254_26034# 6.18e-19
C601 variable_delay_dummy_0.out uio_in[5] 0.11935f
C602 a_25060_23158# ui_in[3] 0.002391f
C603 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.53e-19
C604 variable_delay_short_0.variable_delay_unit_3.in ui_in[2] 3.31e-20
C605 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.53e-19
C606 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward 0.234428f
C607 a_12308_24168# uo_out[1] 6.49e-20
C608 a_24240_11366# ui_in[3] 0.001719f
C609 input_stage_0.fine_delay_unit_1.in uio_in[3] 0.010396f
C610 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.in 7.91e-21
C611 uio_in[4] uio_in[1] 5.22e-19
C612 ui_in[3] ui_in[2] 5.80246f
C613 uio_in[3] uio_in[2] 8.07582f
C614 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_10108_23452# 1.06381f
C615 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_25060_18144# 0.15982f
C616 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12310_39680# 0.014814f
C617 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 uo_out[6] 3.69e-19
C618 uio_oe[1] uio_oe[0] 0.170937f
C619 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[3] 0.014554f
C620 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.010157f
C621 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 5.07283f
C622 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.283838f
C623 a_13254_30598# uo_out[3] 0.188081f
C624 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.283838f
C625 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.871529f
C626 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.003768f
C627 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C628 ui_in[7] uio_in[3] 1.26e-19
C629 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.36e-21
C630 a_12420_33258# uo_out[4] 0.013457f
C631 uio_out[4] uio_out[3] 0.170937f
C632 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 4.28924f
C633 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 uo_out[1] 6.28e-22
C634 a_15322_7112# uio_in[1] 0.003341f
C635 a_9330_14634# VDPWR 1.15434f
C636 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.out 0.172055f
C637 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 3.23832f
C638 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_13254_26034# 0.010872f
C639 VDPWR a_24240_12248# 1.6584f
C640 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.003768f
C641 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_16500_14582# 2.39e-19
C642 VDPWR a_25060_18144# 0.001468f
C643 variable_delay_short_0.out a_16292_8080# 3.3e-19
C644 a_24240_15196# variable_delay_short_0.variable_delay_unit_1.in 7.65e-21
C645 VDPWR a_13254_28694# 6.18e-19
C646 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.in 7.65e-21
C647 uo_out[6] uo_out[5] 1.21073f
C648 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 6.93e-19
C649 a_24240_21092# variable_delay_short_0.variable_delay_unit_3.out 0.493816f
C650 uo_out[7] uo_out[4] 2.26e-21
C651 ui_in[5] uio_in[0] 3e-19
C652 a_12420_33258# a_13254_33258# 0.003413f
C653 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.441213f
C654 a_15680_11634# a_16500_11634# 0.004142f
C655 a_24240_15196# ui_in[7] 0.124274f
C656 a_25060_21092# ui_in[3] 0.002391f
C657 variable_delay_short_0.variable_delay_unit_5.out ui_in[5] 1.07e-20
C658 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_10108_28016# 0.007929f
C659 a_15322_7112# input_stage_0.nand_gate_0.out 3.78e-19
C660 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.499806f
C661 ui_in[5] uio_in[1] 1.46e-19
C662 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.085059f
C663 a_24240_14314# VDPWR 1.6584f
C664 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.in 7.65e-21
C665 variable_delay_short_0.variable_delay_unit_5.out a_24240_26106# 0.505512f
C666 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12310_25988# 0.014814f
C667 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.04313f
C668 uo_out[3] uo_out[2] 2.27264f
C669 a_12420_37822# uo_out[6] 0.013457f
C670 uo_out[4] uo_out[1] 2.26e-21
C671 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_13254_30976# 0.012202f
C672 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.45e-19
C673 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_24240_17262# 0.11539f
C674 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.09966f
C675 a_12308_33296# a_12310_32834# 0.00595f
C676 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_32880# 0.013457f
C677 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.814958f
C678 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.out 0.172055f
C679 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.out 0.085059f
C680 VDPWR a_24240_20210# 1.6584f
C681 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.in 7.65e-21
C682 a_16786_5138# uio_in[5] 0.009499f
C683 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_10108_39426# 0.09966f
C684 VDPWR a_12310_35116# 1.42789f
C685 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en ui_in[3] 0.014554f
C686 a_24790_8314# ui_in[3] 0.024305f
C687 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 8.54e-19
C688 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_24130# 0.504416f
C689 variable_delay_short_0.variable_delay_unit_4.in a_25060_20210# 0.054206f
C690 a_12308_24168# a_13254_24130# 1.02e-19
C691 tdc_0.start_buffer_0.start_buff tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.751615f
C692 variable_delay_short_0.out uio_in[5] 0.075451f
C693 variable_delay_short_0.variable_delay_unit_4.out a_24240_23158# 0.505512f
C694 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.006183f
C695 a_24240_24040# variable_delay_short_0.variable_delay_unit_4.in 7.65e-21
C696 VDPWR uio_in[6] 1.37009f
C697 a_12420_39726# a_13254_39726# 0.003413f
C698 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.006183f
C699 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.15e-21
C700 VDPWR a_24240_17262# 1.6584f
C701 VDPWR variable_delay_short_0.variable_delay_unit_3.in 2.12807f
C702 a_12420_37444# VDPWR 0.497771f
C703 ui_in[4] ui_in[5] 3.94805f
C704 a_25060_24040# ui_in[2] 3.98e-20
C705 VDPWR ui_in[3] 0.206858f
C706 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.out 0.235667f
C707 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 uo_out[6] 6.28e-22
C708 variable_delay_dummy_0.in uio_in[6] 5.32e-19
C709 input_stage_andpwr_0.fine_delay_unit_0.in ua[0] 1.23268f
C710 a_24240_26106# ui_in[4] 0.00352f
C711 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.401225f
C712 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 9.61e-20
C713 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 3.23832f
C714 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12308_31014# 0.162625f
C715 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.138497f
C716 a_16292_6702# uio_in[1] 0.022338f
C717 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.019931f
C718 VDPWR variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 3.87518f
C719 VDPWR a_9330_15794# 1.86061f
C720 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en ui_in[4] 1.11761f
C721 a_12308_35578# a_12420_35540# 0.030083f
C722 VDPWR tdc_0.diff_gen_0.delay_unit_2_5.in_2 3.06042f
C723 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_25060_12248# 0.15982f
C724 variable_delay_dummy_0.variable_delay_unit_1.in a_15680_11634# 0.088132f
C725 ui_in[1] ui_in[0] 6.25329f
C726 uio_in[1] uio_in[5] 3.32e-20
C727 variable_delay_short_0.out variable_delay_dummy_0.out 1.03552f
C728 input_stage_andpwr_0.fine_delay_unit_1.in ui_in[3] 0.020481f
C729 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 9.61e-20
C730 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 2.43248f
C731 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.132512f
C732 a_25060_12248# variable_delay_short_0.in 7.65e-21
C733 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12310_37398# 0.196592f
C734 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.in 0.091118f
C735 a_12420_30598# a_13254_30598# 0.003413f
C736 a_23820_7082# a_24790_6672# 0.53267f
C737 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12310_28270# 0.196592f
C738 a_16292_6702# input_stage_0.nand_gate_0.out 5.26e-20
C739 a_12310_39680# a_12308_37860# 0.005984f
C740 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_25060_26106# 2.39e-19
C741 input_stage_andpwr_0.fine_delay_unit_0.in a_24790_6936# 0.028846f
C742 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.018644f
C743 tdc_0.diff_gen_0.delay_unit_2_3.in_2 a_9330_15794# 0.00105f
C744 a_12420_32880# uo_out[4] 0.492009f
C745 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C746 VDPWR tdc_0.diff_gen_0.delay_unit_2_4.in_2 3.06175f
C747 variable_delay_short_0.variable_delay_unit_4.out a_24240_21092# 0.071074f
C748 input_stage_0.nand_gate_0.out uio_in[5] 0.283562f
C749 variable_delay_dummy_0.variable_delay_unit_1.forward VDPWR 2.28565f
C750 a_24240_23158# a_25060_23158# 0.004142f
C751 VDPWR a_7140_10670# 1.86276f
C752 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.2373f
C753 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.752988f
C754 a_25060_18144# ui_in[5] 6.99e-20
C755 a_15322_8490# uio_in[6] 1.82e-20
C756 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_13254_40104# 0.012202f
C757 uio_oe[6] uio_oe[5] 0.170937f
C758 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_1.in 0.499092f
C759 VDPWR a_12310_28270# 1.42789f
C760 input_stage_andpwr_0.nand_gate_0.out ua[0] 1.24557f
C761 variable_delay_dummy_0.out uio_in[1] 0.001132f
C762 a_9330_15504# a_9330_15794# 0.087529f
C763 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.752988f
C764 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.out 0.493816f
C765 uio_in[7] uio_in[6] 0.073214f
C766 VDPWR tdc_0.diff_gen_0.delay_unit_2_2.in_2 3.0616f
C767 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.04313f
C768 variable_delay_short_0.variable_delay_unit_1.out ui_in[7] 0.224474f
C769 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.953579f
C770 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VDPWR 0.706518f
C771 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 1.24e-19
C772 a_12420_24130# a_13254_24130# 0.003413f
C773 a_12308_24168# VDPWR 1.40782f
C774 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 5.04e-20
C775 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.197073f
C776 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14924# 6.93e-19
C777 a_9330_13764# VDPWR 1.15414f
C778 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.in 0.499092f
C779 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.28924f
C780 a_12420_37444# uo_out[6] 0.492009f
C781 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12310_30552# 0.164402f
C782 a_15322_7112# uio_in[6] 1.82e-20
C783 a_24790_6936# input_stage_andpwr_0.nand_gate_0.out 4.47e-20
C784 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[4] 0.001173f
C785 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.28924f
C786 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_12308_26450# 5.04e-20
C787 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.231672f
C788 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.04313f
C789 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_32880# 0.005542f
C790 rst_n clk 0.031023f
C791 a_24240_20210# ui_in[5] 0.043085f
C792 VDPWR tdc_0.diff_gen_0.delay_unit_2_4.in_1 4.44109f
C793 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.in 0.499092f
C794 a_15680_12516# uio_in[6] 0.001549f
C795 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.231672f
C796 a_24790_8050# ui_in[1] 7.45e-19
C797 a_12310_28270# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 3.45e-19
C798 uo_out[0] uio_in[6] 2.06457f
C799 a_25060_24040# VDPWR 0.001538f
C800 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_23752# 0.013457f
C801 a_12308_24168# a_12310_23706# 0.00595f
C802 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C803 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.start_pos 0.754929f
C804 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 2.43248f
C805 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 7.91e-21
C806 a_9330_15504# tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.001226f
C807 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_4.in 0.499092f
C808 a_24240_26988# ui_in[4] 0.005915f
C809 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.441213f
C810 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12420_30976# 0.003607f
C811 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 uo_out[3] 0.20241f
C812 VDPWR tdc_0.diff_gen_0.delay_unit_2_2.in_1 4.44107f
C813 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[6] 1.53e-22
C814 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.401225f
C815 variable_delay_short_0.variable_delay_unit_3.in ui_in[5] 0.506427f
C816 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_1 0.311186f
C817 a_13254_37444# VDPWR 6.18e-19
C818 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 7.19e-22
C819 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_15680_12516# 0.029284f
C820 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 6.08e-20
C821 a_16500_15464# VDPWR 0.003377f
C822 input_stage_andpwr_0.fine_delay_unit_0.in input_stage_andpwr_0.nand_gate_0.out 0.062321f
C823 variable_delay_short_0.variable_delay_unit_4.in ui_in[6] 0.001632f
C824 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 a_12308_37860# 5.04e-20
C825 ui_in[5] ui_in[3] 0.014973f
C826 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.499806f
C827 variable_delay_short_0.variable_delay_unit_5.in ui_in[4] 0.607531f
C828 a_12310_28270# a_12308_26450# 0.005984f
C829 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_12420_32880# 1.47e-19
C830 a_25060_12248# ui_in[7] 6.99e-20
C831 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.010157f
C832 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 4.53e-19
C833 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_25060_26988# 0.15982f
C834 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq uo_out[5] 0.229249f
C835 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.401225f
C836 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.311186f
C837 variable_delay_short_0.variable_delay_unit_2.out ui_in[7] 0.043504f
C838 a_10108_34862# a_12310_35116# 2.08e-21
C839 a_24240_26106# ui_in[3] 0.001719f
C840 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35540# 0.174293f
C841 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_2 0.667766f
C842 variable_delay_short_0.variable_delay_unit_5.forward a_25060_26106# 0.054206f
C843 VDPWR uo_out[4] 0.587468f
C844 variable_delay_short_0.out uio_in[0] 0.371181f
C845 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en ui_in[3] 0.014554f
C846 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.871529f
C847 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.283838f
C848 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.747722f
C849 a_25060_14314# variable_delay_short_0.variable_delay_unit_1.in 8.82e-20
C850 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en uio_in[6] 0.021622f
C851 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.871529f
C852 a_12310_28270# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.15e-21
C853 variable_delay_short_0.out uio_in[1] 0.030581f
C854 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[4] 0.10528f
C855 a_13254_32880# uo_out[4] 0.188081f
C856 a_24240_23158# VDPWR 1.6584f
C857 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1 0.756572f
C858 a_24240_21092# a_25060_21092# 0.011184f
C859 a_25060_14314# ui_in[7] 0.15982f
C860 a_12308_28732# uo_out[2] 0.014835f
C861 a_25060_23158# variable_delay_short_0.variable_delay_unit_4.in 8.82e-20
C862 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 6.93e-19
C863 a_13254_33258# VDPWR 6.18e-19
C864 input_stage_0.nand_gate_0.out a_16786_5138# 0.355469f
C865 VDPWR a_16500_11634# 0.160518f
C866 a_12420_24130# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.033952f
C867 a_12420_24130# VDPWR 0.497547f
C868 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 3.26e-19
C869 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12310_39680# 0.164402f
C870 uio_in[5] uio_in[6] 5.41755f
C871 a_12308_37860# a_12420_37822# 0.030083f
C872 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.002365f
C873 variable_delay_short_0.variable_delay_unit_4.in ui_in[2] 3.31e-20
C874 a_12420_26034# a_13254_26034# 0.003413f
C875 a_12308_28732# a_12420_28694# 0.030083f
C876 a_9330_14924# VDPWR 1.1544f
C877 uio_in[0] uio_in[1] 6.17178f
C878 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12308_26450# 3.26e-19
C879 a_13254_33258# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.012202f
C880 a_12420_32880# a_12310_32834# 0.030392f
C881 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.756572f
C882 a_24240_11366# a_25060_11366# 0.004142f
C883 a_16500_11634# variable_delay_dummy_0.in 8.82e-20
C884 a_12308_24168# uo_out[0] 0.014835f
C885 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_10108_34862# 0.09966f
C886 tdc_0.start_buffer_0.start_delay variable_delay_short_0.out 6.15e-19
C887 a_25060_11366# ui_in[2] 3.98e-20
C888 ui_in[2] ui_in[0] 0.001501f
C889 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_12310_28270# 3.84e-19
C890 a_23820_8460# ui_in[2] 0.003402f
C891 a_12420_23752# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 1.47e-19
C892 VDPWR tdc_0.vernier_delay_line_0.start_pos 4.78299f
C893 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12420_40104# 0.003607f
C894 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 6.93e-19
C895 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.start_pos 0.283838f
C896 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[5] 0.026424f
C897 a_13254_37444# uo_out[6] 0.188081f
C898 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_1.in 0.087283f
C899 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C900 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_12420_26034# 1.47e-19
C901 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 3.6e-19
C902 a_12420_40104# uo_out[7] 0.013457f
C903 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.forward 0.794183f
C904 variable_delay_dummy_0.out uio_in[6] 0.028463f
C905 input_stage_0.nand_gate_0.out uio_in[1] 1.7e-19
C906 a_24240_21092# VDPWR 1.6584f
C907 variable_delay_short_0.variable_delay_unit_2.in ui_in[7] 0.574722f
C908 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_23752# 0.005542f
C909 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_10108_25734# 0.192064f
C910 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12308_37860# 3.26e-19
C911 uio_oe[0] uio_out[7] 0.170937f
C912 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57489f
C913 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.2373f
C914 ua[0] uio_in[6] 0.243341f
C915 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 4.28924f
C916 ui_in[4] uio_in[0] 1.15e-19
C917 variable_delay_short_0.variable_delay_unit_5.out ui_in[4] 0.047464f
C918 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12420_30598# 0.035356f
C919 uo_out[6] uo_out[4] 1.58e-19
C920 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.6e-19
C921 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 1.17e-19
C922 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 a_12308_35578# 5.04e-20
C923 a_13254_35540# uo_out[5] 0.005542f
C924 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.162625f
C925 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 VDPWR 5.07283f
C926 uio_out[3] uio_out[2] 0.170937f
C927 a_24240_26988# ui_in[3] 0.001719f
C928 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12308_40142# 0.162625f
C929 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.out 0.12022f
C930 a_16500_11634# uio_in[4] 6.61e-20
C931 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_25060_24040# 0.15982f
C932 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.019931f
C933 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.138497f
C934 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12310_23706# 0.196592f
C935 VDPWR variable_delay_dummy_0.variable_delay_unit_1.in 3.21199f
C936 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 a_12420_37444# 1.47e-19
C937 a_12308_40142# uo_out[7] 0.01561f
C938 a_9330_14634# variable_delay_short_0.out 2.11e-19
C939 variable_delay_short_0.out a_24240_12248# 0.493816f
C940 uo_out[3] uo_out[1] 1.56e-19
C941 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.138497f
C942 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 5.04e-20
C943 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 7.91e-21
C944 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 uo_out[3] 1.35e-20
C945 tdc_0.start_buffer_0.start_buff a_9330_14054# 1.66e-19
C946 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12310_35116# 0.014814f
C947 variable_delay_short_0.variable_delay_unit_5.in ui_in[3] 0.02f
C948 a_24240_15196# variable_delay_short_0.variable_delay_unit_1.out 0.493816f
C949 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 9.61e-20
C950 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_24240_11366# 0.11539f
C951 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.in 0.08442f
C952 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en ui_in[2] 6.97e-19
C953 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.018644f
C954 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 3.6e-19
C955 a_12420_28694# uo_out[2] 0.013457f
C956 a_24790_8050# ui_in[2] 0.023539f
C957 a_23820_8460# a_24790_8314# 0.019821f
C958 a_24240_11366# variable_delay_short_0.in 8.82e-20
C959 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.002365f
C960 variable_delay_dummy_0.out a_7140_10670# 0.087271f
C961 variable_delay_short_0.in ui_in[2] 1.86e-20
C962 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.003768f
C963 a_24240_12248# uio_in[0] 0.124274f
C964 a_12310_37398# a_12308_35578# 0.005984f
C965 variable_delay_short_0.variable_delay_unit_4.in VDPWR 2.12807f
C966 a_12420_24130# uo_out[0] 0.013457f
C967 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_16500_15464# 0.15982f
C968 a_12310_32834# VDPWR 1.42789f
C969 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq uo_out[1] 0.229249f
C970 input_stage_andpwr_0.fine_delay_unit_0.in uio_in[6] 3.47e-19
C971 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_12310_28270# 4.55e-19
C972 VDPWR a_25060_11366# 6.98e-19
C973 VDPWR ui_in[0] 4.76e-19
C974 a_12420_23752# VDPWR 0.497771f
C975 a_23820_8460# VDPWR 1.25074f
C976 a_12420_23752# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.003664f
C977 a_10108_37144# a_12310_37398# 2.08e-21
C978 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12308_26450# 2.36e-21
C979 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37822# 0.174293f
C980 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28694# 0.174293f
C981 a_16786_5138# uio_in[6] 0.010606f
C982 a_10108_28016# a_12310_28270# 2.08e-21
C983 a_23820_7082# ui_in[1] 0.010812f
C984 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_24240_23158# 0.11539f
C985 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.164402f
C986 ui_in[6] uio_in[2] 1.69e-19
C987 a_12310_32834# a_13254_32880# 1.02e-19
C988 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.231672f
C989 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C990 variable_delay_short_0.out uio_in[6] 0.02732f
C991 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.002141f
C992 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.forward 0.794183f
C993 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12308_28732# 7.19e-22
C994 variable_delay_dummy_0.variable_delay_unit_1.in uio_in[4] 4.58e-20
C995 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.36e-21
C996 a_12420_23752# a_12310_23706# 0.030392f
C997 a_23820_8460# input_stage_andpwr_0.fine_delay_unit_1.in 0.254332f
C998 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_10108_25734# 0.007929f
C999 ui_in[6] ui_in[7] 7.62803f
C1000 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.747722f
C1001 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12420_39726# 0.035356f
C1002 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.out 0.071074f
C1003 variable_delay_short_0.out ui_in[3] 0.06888f
C1004 a_12420_33258# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.003607f
C1005 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2 0.04313f
C1006 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12308_35578# 3.26e-19
C1007 a_12420_39726# uo_out[7] 0.492009f
C1008 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 uo_out[0] 0.20241f
C1009 a_12308_31014# VDPWR 1.40782f
C1010 input_stage_andpwr_0.nand_gate_0.out uio_in[6] 0.052822f
C1011 variable_delay_short_0.out variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 2.24e-20
C1012 a_24790_8314# a_24790_8050# 0.556904f
C1013 variable_delay_dummy_0.variable_delay_unit_1.forward a_16500_14582# 0.054206f
C1014 a_24240_21092# ui_in[5] 0.124669f
C1015 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.441213f
C1016 variable_delay_dummy_0.variable_delay_unit_1.out a_16500_12516# 0.070146f
C1017 a_24790_8314# variable_delay_short_0.in 7.3e-20
C1018 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_10108_37144# 0.09966f
C1019 variable_delay_dummy_0.variable_delay_unit_1.in a_15680_12516# 0.020173f
C1020 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_13254_30598# 0.010872f
C1021 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 6.08e-20
C1022 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 uo_out[3] 3.69e-19
C1023 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_10108_28016# 0.09966f
C1024 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 3.26e-19
C1025 uio_in[0] ui_in[3] 0.014973f
C1026 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_25060_20210# 2.39e-19
C1027 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 a_12420_35162# 1.47e-19
C1028 a_12310_35116# uo_out[5] 0.098308f
C1029 a_16500_11634# uio_in[5] 0.002787f
C1030 variable_delay_short_0.variable_delay_unit_5.out ui_in[3] 0.040959f
C1031 variable_delay_short_0.variable_delay_unit_1.in a_24240_11366# 0.088132f
C1032 variable_delay_short_0.variable_delay_unit_1.in ui_in[2] 3.31e-20
C1033 VDPWR variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 2.78173f
C1034 uio_oe[5] uio_oe[4] 0.170937f
C1035 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.in 0.09141f
C1036 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 9.61e-20
C1037 input_stage_0.nand_gate_0.out uio_in[6] 0.054416f
C1038 a_12420_30598# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 1.47e-19
C1039 VDPWR variable_delay_short_0.in 1.34358f
C1040 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.53e-19
C1041 ui_in[7] ui_in[2] 7.13e-19
C1042 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.out 0.12029f
C1043 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_5.in_2 0.401225f
C1044 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[7] 1.09349f
C1045 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.667766f
C1046 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1047 a_12420_28316# uo_out[2] 0.492009f
C1048 a_13254_26412# uo_out[1] 0.005542f
C1049 a_24790_6672# ui_in[1] 0.00799f
C1050 input_stage_andpwr_0.fine_delay_unit_1.in a_24790_8050# 0.244525f
C1051 a_24240_18144# variable_delay_short_0.variable_delay_unit_2.out 0.493816f
C1052 variable_delay_dummy_0.out a_16500_11634# 0.222585f
C1053 a_25060_15196# ui_in[3] 0.002391f
C1054 input_stage_andpwr_0.fine_delay_unit_1.in variable_delay_short_0.in 0.002949f
C1055 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.100263f
C1056 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 uo_out[6] 0.20241f
C1057 clk ena 0.031023f
C1058 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[5] 0.10528f
C1059 ui_in[4] ui_in[3] 2.58276f
C1060 variable_delay_short_0.variable_delay_unit_4.in ui_in[5] 0.586739f
C1061 a_12420_23752# uo_out[0] 0.492009f
C1062 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_13254_35540# 0.012202f
C1063 a_9330_13764# variable_delay_short_0.out 0.076613f
C1064 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.007929f
C1065 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.in 0.020173f
C1066 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.in 0.09141f
C1067 a_12420_40104# VDPWR 0.497547f
C1068 a_9330_14344# a_9330_14054# 0.083149f
C1069 a_13254_23752# VDPWR 6.18e-19
C1070 a_24240_23158# variable_delay_short_0.variable_delay_unit_5.in 0.088132f
C1071 variable_delay_dummy_0.variable_delay_unit_1.out a_15680_14582# 0.505512f
C1072 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12310_37398# 0.014814f
C1073 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12310_28270# 0.014814f
C1074 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.in 0.09141f
C1075 variable_delay_dummy_0.in a_16292_8344# 7.3e-20
C1076 a_25060_26106# ui_in[2] 3.98e-20
C1077 a_12420_30976# VDPWR 0.497547f
C1078 VDPWR uo_out[3] 0.587468f
C1079 variable_delay_dummy_0.variable_delay_unit_1.in uio_in[5] 0.019965f
C1080 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.99e-19
C1081 a_12310_23706# a_13254_23752# 1.02e-19
C1082 a_9330_15214# VDPWR 1.15434f
C1083 tdc_0.start_buffer_0.start_delay a_7140_10670# 7.1e-20
C1084 variable_delay_short_0.variable_delay_unit_1.out a_25060_12248# 0.070146f
C1085 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_13254_39726# 0.010872f
C1086 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.out 0.071795f
C1087 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[3] 6.28e-22
C1088 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.953579f
C1089 a_12308_40142# VDPWR 1.40742f
C1090 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.953579f
C1091 a_13254_39726# uo_out[7] 0.188251f
C1092 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en ui_in[7] 1.5e-19
C1093 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1 0.001356f
C1094 a_12420_32880# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.035356f
C1095 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.6e-19
C1096 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12308_35578# 0.162625f
C1097 a_25060_24040# variable_delay_short_0.variable_delay_unit_5.out 0.070146f
C1098 variable_delay_short_0.variable_delay_unit_3.out a_24240_18144# 0.071074f
C1099 a_24240_12248# ui_in[3] 0.001719f
C1100 VDPWR input_stage_0.fine_delay_unit_1.in 1.33446f
C1101 VDPWR uio_in[2] 0.005628f
C1102 VDPWR variable_delay_short_0.variable_delay_unit_1.in 2.13093f
C1103 a_25060_18144# ui_in[3] 0.002391f
C1104 a_9330_14634# a_9330_15794# 2.78e-19
C1105 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.706518f
C1106 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.out 0.235655f
C1107 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.231672f
C1108 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.231672f
C1109 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[4] 1.53e-22
C1110 tdc_0.start_buffer_0.start_delay a_9330_13764# 1.56e-19
C1111 variable_delay_short_0.variable_delay_unit_1.out a_25060_14314# 0.222585f
C1112 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.006183f
C1113 a_24240_18144# variable_delay_short_0.variable_delay_unit_2.in 7.65e-21
C1114 ui_in[6] uio_in[3] 9.55e-20
C1115 a_15322_8490# a_16292_8344# 0.019821f
C1116 a_12420_35162# a_13254_35162# 0.003413f
C1117 VDPWR ui_in[7] 1.41097f
C1118 variable_delay_dummy_0.in input_stage_0.fine_delay_unit_1.in 0.002924f
C1119 a_9330_15504# a_9330_15214# 0.083149f
C1120 a_16292_8344# uio_in[4] 0.024305f
C1121 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.018644f
C1122 variable_delay_dummy_0.in uio_in[2] 1.05e-20
C1123 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.085059f
C1124 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[3] 3.5e-20
C1125 input_stage_0.fine_delay_unit_0.in VDPWR 1.53841f
C1126 VDPWR tdc_0.diff_gen_0.delay_unit_2_1.in_1 4.44048f
C1127 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 2.59e-20
C1128 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.in 8.82e-20
C1129 a_24240_14314# ui_in[3] 0.001719f
C1130 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12310_25988# 6.08e-20
C1131 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30976# 0.504416f
C1132 a_12308_31014# a_13254_30976# 1.02e-19
C1133 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq uo_out[3] 0.229249f
C1134 VDPWR a_16500_12516# 0.003447f
C1135 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en ui_in[6] 4.42e-19
C1136 a_24240_20210# ui_in[3] 0.001719f
C1137 a_25060_24040# ui_in[4] 0.001909f
C1138 a_9330_14924# variable_delay_short_0.out 8.85e-20
C1139 a_12310_25988# uo_out[1] 0.098308f
C1140 a_24240_15196# ui_in[6] 6.99e-20
C1141 a_13254_28316# uo_out[2] 0.188081f
C1142 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.132512f
C1143 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.vernier_delay_line_0.start_pos 0.400636f
C1144 variable_delay_short_0.variable_delay_unit_3.in a_24240_17262# 0.088132f
C1145 variable_delay_short_0.variable_delay_unit_1.out ui_in[1] 0.001119f
C1146 a_16500_12516# variable_delay_dummy_0.in 7.65e-21
C1147 uo_out[6] uo_out[3] 2.26e-21
C1148 uo_out[5] uo_out[4] 1.5647f
C1149 a_24240_17262# ui_in[3] 0.001719f
C1150 variable_delay_short_0.variable_delay_unit_3.in ui_in[3] 0.02f
C1151 rst_n ui_in[0] 0.031023f
C1152 a_15322_8490# input_stage_0.fine_delay_unit_1.in 0.254332f
C1153 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12310_35116# 0.164402f
C1154 a_13254_23752# uo_out[0] 0.188081f
C1155 a_25060_26988# ui_in[2] 3.98e-20
C1156 VDPWR a_25060_26106# 0.160518f
C1157 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 1.24e-19
C1158 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 0.002141f
C1159 ua[0] ui_in[0] 1.96e-19
C1160 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[6] 0.013186f
C1161 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in 0.235667f
C1162 input_stage_0.fine_delay_unit_1.in uio_in[4] 0.020481f
C1163 a_12420_39726# VDPWR 0.497771f
C1164 a_9330_15504# tdc_0.diff_gen_0.delay_unit_2_1.in_1 8.59e-20
C1165 uio_in[4] uio_in[2] 0.01853f
C1166 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_5.in 0.087283f
C1167 a_16500_14582# variable_delay_dummy_0.variable_delay_unit_1.in 8.82e-20
C1168 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[6] 2.92e-19
C1169 uo_out[3] uo_out[0] 2.26e-21
C1170 uo_out[2] uo_out[1] 2.62662f
C1171 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1172 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.100263f
C1173 ui_in[7] uio_in[4] 3.77e-20
C1174 a_15322_7112# a_16292_6966# 0.019821f
C1175 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1176 a_12420_40104# a_13254_40104# 0.003413f
C1177 a_16292_8344# a_16292_8080# 0.556904f
C1178 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.36e-21
C1179 uio_out[2] uio_out[1] 0.170937f
C1180 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12420_35540# 0.003607f
C1181 a_15322_7112# input_stage_0.fine_delay_unit_1.in 0.130264f
C1182 a_12420_30598# VDPWR 0.497771f
C1183 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en ui_in[2] 6.97e-19
C1184 VDPWR tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.57093f
C1185 VDPWR a_12308_35578# 1.40782f
C1186 a_24790_6936# ui_in[0] 0.022567f
C1187 a_15322_7112# uio_in[2] 0.010812f
C1188 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.vernier_delay_line_0.start_pos 0.728719f
C1189 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.001356f
C1190 a_24240_23158# ui_in[4] 0.046238f
C1191 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.499806f
C1192 variable_delay_dummy_0.variable_delay_unit_1.forward uio_in[6] 0.03353f
C1193 VDPWR a_13254_26412# 6.18e-19
C1194 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.003768f
C1195 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_13254_37822# 0.012202f
C1196 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.231672f
C1197 a_15680_14582# VDPWR 1.70112f
C1198 a_16500_12516# uio_in[4] 6.61e-20
C1199 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.28924f
C1200 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_13254_28694# 0.012202f
C1201 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.45e-19
C1202 a_13254_32880# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.010872f
C1203 variable_delay_short_0.variable_delay_unit_2.out a_25060_17262# 0.222585f
C1204 a_23820_7082# VDPWR 1.25313f
C1205 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12310_35116# 6.08e-20
C1206 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_24240_15196# 0.029284f
C1207 a_24240_18144# ui_in[6] 0.124274f
C1208 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out 0.071795f
C1209 variable_delay_short_0.variable_delay_unit_2.out ui_in[1] 0.001119f
C1210 a_15322_7112# input_stage_0.fine_delay_unit_0.in 0.254311f
C1211 ui_in[5] uio_in[2] 9.52e-20
C1212 a_12308_40142# a_13254_40104# 1.02e-19
C1213 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12420_40104# 0.504416f
C1214 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.start_buffer_0.start_buff 0.311237f
C1215 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2 0.04313f
C1216 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 7.91e-21
C1217 a_12420_30976# a_13254_30976# 0.003413f
C1218 a_13254_30976# uo_out[3] 0.005542f
C1219 input_stage_andpwr_0.fine_delay_unit_0.in ui_in[0] 0.009426f
C1220 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.59e-20
C1221 input_stage_andpwr_0.fine_delay_unit_1.in a_23820_7082# 0.130264f
C1222 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_2.in 0.499092f
C1223 input_stage_0.fine_delay_unit_1.in a_16292_8080# 0.244525f
C1224 ui_in[5] ui_in[7] 0.00231f
C1225 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 uo_out[4] 3.69e-19
C1226 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[2] 6.97e-19
C1227 a_16292_8344# uio_in[5] 0.001923f
C1228 a_16292_8080# uio_in[2] 0.001529f
C1229 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.start_neg 0.626611f
C1230 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_25060_21092# 0.15982f
C1231 a_15680_12516# a_16500_12516# 0.011184f
C1232 tdc_0.diff_gen_0.delay_unit_2_2.in_2 a_9330_15794# 0.001232f
C1233 variable_delay_short_0.out a_25060_11366# 0.222585f
C1234 variable_delay_short_0.variable_delay_unit_3.out a_25060_20210# 0.222585f
C1235 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12308_37860# 0.162625f
C1236 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30598# 0.013457f
C1237 a_12308_31014# a_12310_30552# 0.00595f
C1238 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12308_28732# 0.162625f
C1239 a_23820_8460# variable_delay_short_0.out 0.00491f
C1240 a_24240_21092# ui_in[4] 6.99e-20
C1241 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1242 a_25060_14314# variable_delay_short_0.variable_delay_unit_2.in 0.054206f
C1243 input_stage_0.fine_delay_unit_0.in a_16292_8080# 1.39e-20
C1244 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.100263f
C1245 VDPWR a_25060_26988# 0.003377f
C1246 variable_delay_short_0.variable_delay_unit_1.out ui_in[6] 2.67e-19
C1247 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C1248 a_25060_24040# ui_in[3] 0.002391f
C1249 a_16292_6966# a_16292_6702# 0.556904f
C1250 a_9330_14924# a_9330_14634# 0.083149f
C1251 VDPWR uio_in[3] 0.001248f
C1252 variable_delay_dummy_0.out a_16292_8344# 5.64e-19
C1253 a_16500_15464# uio_in[6] 0.002068f
C1254 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_1 0.311186f
C1255 a_12420_37444# a_13254_37444# 0.003413f
C1256 a_16292_6702# input_stage_0.fine_delay_unit_1.in 7.4e-19
C1257 VDPWR a_12308_28732# 1.40782f
C1258 a_25060_11366# uio_in[0] 0.15982f
C1259 input_stage_andpwr_0.nand_gate_0.out ui_in[0] 1.7e-19
C1260 a_16292_6966# uio_in[5] 2.26e-20
C1261 a_12420_28316# a_13254_28316# 0.003413f
C1262 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.018644f
C1263 a_16292_6702# uio_in[2] 0.00799f
C1264 a_12308_26450# a_13254_26412# 1.02e-19
C1265 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26412# 0.504416f
C1266 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.018644f
C1267 a_23820_8460# uio_in[0] 1.26e-19
C1268 variable_delay_short_0.variable_delay_unit_3.out ui_in[1] 0.001119f
C1269 a_12308_35578# uo_out[6] 6.49e-20
C1270 a_12308_33296# a_12420_33258# 0.030083f
C1271 input_stage_0.fine_delay_unit_1.in uio_in[5] 0.011377f
C1272 variable_delay_dummy_0.in uio_in[3] 5.31e-20
C1273 variable_delay_short_0.variable_delay_unit_5.forward ui_in[6] 0.001598f
C1274 a_13254_39726# VDPWR 6.18e-19
C1275 uio_in[2] uio_in[5] 1.37e-20
C1276 VDPWR a_12420_35540# 0.497547f
C1277 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en VDPWR 2.77611f
C1278 tdc_0.diff_gen_0.delay_unit_2_2.in_1 a_9330_15794# 4.02e-19
C1279 a_25060_17262# variable_delay_short_0.variable_delay_unit_2.in 8.82e-20
C1280 a_24790_6672# VDPWR 5.43e-20
C1281 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14054# 8.73e-19
C1282 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.2373f
C1283 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_2 0.667766f
C1284 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_13254_26412# 0.012202f
C1285 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.010157f
C1286 a_24240_26106# a_25060_26106# 0.004142f
C1287 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12308_31014# 0.197073f
C1288 a_24240_15196# VDPWR 1.6584f
C1289 input_stage_0.fine_delay_unit_0.in a_16292_6702# 0.244525f
C1290 a_24790_8050# input_stage_andpwr_0.fine_delay_unit_0.in 1.39e-20
C1291 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.499806f
C1292 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12420_35162# 0.035356f
C1293 a_13254_30598# VDPWR 6.18e-19
C1294 input_stage_0.fine_delay_unit_0.in uio_in[5] 0.042742f
C1295 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 2.36e-21
C1296 input_stage_andpwr_0.fine_delay_unit_1.in a_24790_6672# 7.4e-19
C1297 variable_delay_short_0.variable_delay_unit_4.in ui_in[4] 0.507197f
C1298 variable_delay_dummy_0.out input_stage_0.fine_delay_unit_1.in 0.024958f
C1299 variable_delay_short_0.variable_delay_unit_1.out ui_in[2] 0.002549f
C1300 VDPWR a_12310_25988# 1.42789f
C1301 uio_oe[4] uio_oe[3] 0.170937f
C1302 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12310_37398# 0.164402f
C1303 variable_delay_dummy_0.out uio_in[2] 0.001744f
C1304 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.120255f
C1305 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1306 tdc_0.start_buffer_0.start_buff VDPWR 7.34803f
C1307 a_16500_12516# uio_in[5] 0.002787f
C1308 a_24240_23158# ui_in[3] 0.001719f
C1309 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12310_28270# 0.164402f
C1310 a_24790_8050# variable_delay_short_0.out 6.1e-19
C1311 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.499806f
C1312 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.953579f
C1313 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[4] 6.28e-22
C1314 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.out 0.12029f
C1315 variable_delay_short_0.variable_delay_unit_2.out ui_in[6] 0.224474f
C1316 variable_delay_short_0.out variable_delay_short_0.in 0.599483f
C1317 VDPWR tdc_0.vernier_delay_line_0.start_neg 3.22778f
C1318 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VDPWR 0.706518f
C1319 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.start_neg 0.019727f
C1320 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.007279f
C1321 a_15322_8490# uio_in[3] 0.003646f
C1322 VDPWR variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 3.86957f
C1323 uio_in[4] uio_in[3] 9.04698f
C1324 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 uo_out[2] 0.20241f
C1325 a_25284_5108# VDPWR 0.009499f
C1326 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.667766f
C1327 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_24240_18144# 0.029284f
C1328 variable_delay_short_0.variable_delay_unit_5.forward ui_in[2] 1.68e-20
C1329 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12420_39726# 0.013457f
C1330 a_12308_40142# a_12310_39680# 0.00595f
C1331 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_16500_11634# 2.39e-19
C1332 a_12310_30552# uo_out[3] 0.098308f
C1333 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12420_37822# 0.003607f
C1334 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en uio_in[0] 1.09349f
C1335 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_10108_32580# 0.192064f
C1336 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12420_28694# 0.003607f
C1337 a_16500_12516# variable_delay_dummy_0.out 0.172055f
C1338 VDPWR uo_out[2] 0.587468f
C1339 variable_delay_short_0.in uio_in[0] 0.26219f
C1340 a_9330_14924# a_9330_15794# 4.98e-19
C1341 a_24240_24040# variable_delay_short_0.variable_delay_unit_4.out 0.493816f
C1342 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12310_25988# 0.196592f
C1343 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_15680_14582# 0.11539f
C1344 VDPWR a_24240_18144# 1.6584f
C1345 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.001356f
C1346 variable_delay_short_0.out a_16292_8344# 2.5e-19
C1347 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30598# 0.005542f
C1348 VDPWR a_12420_28694# 0.497547f
C1349 a_12420_26412# a_13254_26412# 0.003413f
C1350 a_24240_21092# variable_delay_short_0.variable_delay_unit_3.in 7.65e-21
C1351 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq uo_out[4] 0.229249f
C1352 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out 0.071795f
C1353 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 4.55e-19
C1354 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14344# 0.001157f
C1355 a_25060_12248# ui_in[2] 3.98e-20
C1356 variable_delay_short_0.variable_delay_unit_4.out ui_in[1] 0.001119f
C1357 a_24240_21092# ui_in[3] 0.001719f
C1358 variable_delay_short_0.variable_delay_unit_2.out ui_in[2] 0.002549f
C1359 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.747722f
C1360 a_25060_17262# ui_in[6] 0.15982f
C1361 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 6.79e-20
C1362 variable_delay_short_0.variable_delay_unit_3.out ui_in[6] 0.043504f
C1363 a_9330_14054# VDPWR 1.1544f
C1364 variable_delay_dummy_0.variable_delay_unit_1.in uio_in[6] 0.018232f
C1365 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 1.17e-19
C1366 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26034# 0.013457f
C1367 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.085059f
C1368 a_12308_26450# a_12310_25988# 0.00595f
C1369 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002141f
C1370 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[3] 0.10528f
C1371 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12420_30976# 0.033952f
C1372 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[7] 1.53e-22
C1373 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.2373f
C1374 a_10108_32580# a_12310_32834# 2.08e-21
C1375 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_33258# 0.174293f
C1376 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 7.19e-22
C1377 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.out 0.493816f
C1378 a_16292_8080# uio_in[3] 0.023966f
C1379 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 VDPWR 5.07283f
C1380 VDPWR a_12420_35162# 0.497771f
C1381 variable_delay_short_0.variable_delay_unit_2.in ui_in[6] 0.50637f
C1382 variable_delay_short_0.variable_delay_unit_4.in a_24240_20210# 0.088132f
C1383 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en ui_in[5] 1.10207f
C1384 a_12308_24168# a_12420_24130# 0.030083f
C1385 a_25060_14314# ui_in[2] 3.98e-20
C1386 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.192064f
C1387 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 uo_out[7] 0.203149f
C1388 variable_delay_short_0.out input_stage_0.fine_delay_unit_1.in 0.008066f
C1389 a_25060_26106# variable_delay_short_0.variable_delay_unit_5.in 8.82e-20
C1390 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_12310_25988# 0.164402f
C1391 variable_delay_short_0.out uio_in[2] 0.022033f
C1392 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.814958f
C1393 variable_delay_short_0.variable_delay_unit_1.out VDPWR 1.34424f
C1394 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq uo_out[6] 0.229249f
C1395 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in 0.235655f
C1396 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.2373f
C1397 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.003768f
C1398 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1399 a_12420_39726# a_12310_39680# 0.030392f
C1400 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_25060_14314# 2.39e-19
C1401 a_25060_20210# ui_in[2] 3.98e-20
C1402 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_13254_35162# 0.010872f
C1403 a_13254_37822# VDPWR 6.18e-19
C1404 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.002365f
C1405 a_12308_26450# uo_out[2] 6.49e-20
C1406 variable_delay_short_0.out ui_in[7] 2.67e-19
C1407 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.in 0.087283f
C1408 VDPWR variable_delay_short_0.variable_delay_unit_5.forward 2.28561f
C1409 a_23820_7082# ua[0] 0.002135f
C1410 variable_delay_short_0.variable_delay_unit_4.in ui_in[3] 0.02f
C1411 tdc_0.diff_gen_0.delay_unit_2_1.in_1 variable_delay_short_0.out 7.3e-20
C1412 a_25060_17262# ui_in[2] 3.98e-20
C1413 a_16292_6966# uio_in[1] 0.022988f
C1414 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_10108_30298# 1.06381f
C1415 uo_out[5] uo_out[3] 1.56e-19
C1416 variable_delay_short_0.variable_delay_unit_1.in uio_in[0] 0.574722f
C1417 a_12310_37398# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 3.45e-19
C1418 variable_delay_short_0.variable_delay_unit_3.out ui_in[2] 0.002549f
C1419 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_24240_12248# 0.029284f
C1420 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.in 0.087283f
C1421 uio_out[6] uio_out[5] 0.170937f
C1422 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 uo_out[2] 1.53e-22
C1423 a_25060_11366# ui_in[3] 0.002391f
C1424 ui_in[3] ui_in[0] 2.87e-19
C1425 uio_in[3] uio_in[5] 0.001464f
C1426 ui_in[2] ui_in[1] 5.7665f
C1427 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[5] 7.3e-19
C1428 uio_in[2] uio_in[1] 9.35827f
C1429 ui_in[7] uio_in[0] 9.98875f
C1430 a_23820_8460# ui_in[3] 0.010812f
C1431 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12308_24168# 0.162625f
C1432 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.12029f
C1433 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 a_10108_37144# 0.192064f
C1434 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_13254_39726# 0.005542f
C1435 a_24240_12248# variable_delay_short_0.in 7.65e-21
C1436 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12420_37444# 0.035356f
C1437 a_12420_30598# a_12310_30552# 0.030392f
C1438 uo_out[2] uo_out[0] 1.56e-19
C1439 a_23820_7082# a_24790_6936# 0.019821f
C1440 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_24240_26106# 0.11539f
C1441 a_16292_6966# input_stage_0.nand_gate_0.out 4.47e-20
C1442 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12420_28316# 0.035356f
C1443 variable_delay_short_0.variable_delay_unit_2.in ui_in[2] 3.31e-20
C1444 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 8.54e-19
C1445 ui_in[7] uio_in[1] 5.13e-19
C1446 a_13254_33258# uo_out[4] 0.005542f
C1447 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.59e-20
C1448 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.100263f
C1449 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.in 0.814958f
C1450 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 0.002365f
C1451 a_9330_14344# VDPWR 1.1544f
C1452 input_stage_0.nand_gate_0.out uio_in[2] 6.37e-19
C1453 input_stage_0.fine_delay_unit_0.in uio_in[1] 0.009426f
C1454 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.6e-19
C1455 VDPWR a_25060_12248# 0.001468f
C1456 VDPWR variable_delay_short_0.variable_delay_unit_2.out 1.34424f
C1457 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12420_40104# 0.033952f
C1458 a_24240_18144# ui_in[5] 6.99e-20
C1459 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.in 7.65e-21
C1460 VDPWR a_12420_28316# 0.497771f
C1461 variable_delay_dummy_0.out uio_in[3] 0.002875f
C1462 a_24240_26988# a_25060_26988# 0.011184f
C1463 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 uo_out[2] 1.35e-20
C1464 a_15680_14582# a_16500_14582# 0.004142f
C1465 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.out 0.172055f
C1466 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 6.79e-20
C1467 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.747722f
C1468 uio_out[1] uio_out[0] 0.170937f
C1469 a_25060_15196# ui_in[7] 0.001909f
C1470 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C1471 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 VDPWR 3.23832f
C1472 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_12308_28732# 5.04e-20
C1473 a_23820_7082# input_stage_andpwr_0.fine_delay_unit_0.in 0.254311f
C1474 a_12308_33296# VDPWR 1.40782f
C1475 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out 0.062023f
C1476 ui_in[4] ui_in[7] 0.002007f
C1477 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.09966f
C1478 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.007929f
C1479 tdc_0.start_buffer_0.start_delay tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.401491f
C1480 a_25060_14314# VDPWR 6.98e-19
C1481 variable_delay_short_0.variable_delay_unit_5.out a_25060_26106# 0.222585f
C1482 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26034# 0.005542f
C1483 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.in 7.65e-21
C1484 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12420_30598# 0.003664f
C1485 a_13254_37822# uo_out[6] 0.005542f
C1486 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.747722f
C1487 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 9.61e-20
C1488 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 6.79e-20
C1489 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.197073f
C1490 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_25060_17262# 2.39e-19
C1491 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12310_32834# 0.014814f
C1492 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.085059f
C1493 VDPWR a_25060_20210# 6.98e-19
C1494 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12308_40142# 0.197073f
C1495 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en ui_in[3] 0.014554f
C1496 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.in 7.65e-21
C1497 VDPWR a_13254_35162# 6.18e-19
C1498 a_24790_8314# ui_in[1] 4.3e-19
C1499 a_24790_8050# ui_in[3] 0.00799f
C1500 a_24240_24040# VDPWR 1.65847f
C1501 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_24130# 0.174293f
C1502 a_10108_23452# a_12310_23706# 2.08e-21
C1503 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 8.54e-19
C1504 variable_delay_short_0.in ui_in[3] 0.052959f
C1505 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 uo_out[4] 1.35e-20
C1506 uio_out[0] uo_out[7] 0.170937f
C1507 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.in 7.65e-21
C1508 variable_delay_short_0.variable_delay_unit_4.out a_25060_23158# 0.222585f
C1509 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 8.54e-19
C1510 a_12310_39680# a_13254_39726# 1.02e-19
C1511 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.in 7.91e-21
C1512 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.in 0.09141f
C1513 VDPWR a_25060_17262# 6.98e-19
C1514 tdc_0.start_buffer_0.start_buff variable_delay_dummy_0.out 5.26e-19
C1515 a_12310_37398# VDPWR 1.42789f
C1516 VDPWR variable_delay_short_0.variable_delay_unit_3.out 1.34424f
C1517 variable_delay_short_0.variable_delay_unit_1.in a_24240_12248# 0.020173f
C1518 a_12310_30552# a_12308_28732# 0.005984f
C1519 variable_delay_short_0.variable_delay_unit_4.out ui_in[2] 0.002549f
C1520 a_23820_7082# input_stage_andpwr_0.nand_gate_0.out 3.78e-19
C1521 a_15680_15464# VDPWR 1.78268f
C1522 a_24790_6936# a_24790_6672# 0.556904f
C1523 VDPWR ui_in[1] 0.002882f
C1524 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12420_24130# 0.003607f
C1525 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 a_10108_37144# 0.007929f
C1526 variable_delay_short_0.variable_delay_unit_5.forward ui_in[5] 0.003308f
C1527 a_24240_12248# ui_in[7] 6.99e-20
C1528 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.132512f
C1529 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_24240_26988# 0.029284f
C1530 a_12308_35578# uo_out[5] 0.014835f
C1531 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.953579f
C1532 ui_in[6] ui_in[2] 7.13e-19
C1533 VDPWR variable_delay_short_0.variable_delay_unit_2.in 2.12807f
C1534 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 a_10108_34862# 0.192064f
C1535 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35540# 0.504416f
C1536 a_12308_35578# a_13254_35540# 1.02e-19
C1537 a_25284_5108# ua[0] 7.57e-19
C1538 variable_delay_dummy_0.variable_delay_unit_1.in a_16500_11634# 0.054206f
C1539 variable_delay_short_0.variable_delay_unit_5.forward a_24240_26106# 0.088132f
C1540 ua[1] VGND 0.146962f
C1541 ua[2] VGND 0.146962f
C1542 ua[3] VGND 0.146962f
C1543 ua[4] VGND 0.146962f
C1544 ua[5] VGND 0.146962f
C1545 ua[6] VGND 0.146962f
C1546 ua[7] VGND 0.146962f
C1547 ena VGND 0.070385f
C1548 clk VGND 0.042875f
C1549 rst_n VGND 0.042875f
C1550 uio_in[7] VGND 0.071255f
C1551 uio_out[0] VGND 0.136988f
C1552 uio_out[1] VGND 0.136988f
C1553 uio_out[2] VGND 0.137343f
C1554 uio_out[3] VGND 0.137343f
C1555 uio_out[4] VGND 0.137343f
C1556 uio_out[5] VGND 0.137343f
C1557 uio_out[6] VGND 0.137343f
C1558 uio_out[7] VGND 0.137343f
C1559 uio_oe[0] VGND 0.137343f
C1560 uio_oe[1] VGND 0.137343f
C1561 uio_oe[2] VGND 0.137343f
C1562 uio_oe[3] VGND 0.137339f
C1563 uio_oe[4] VGND 0.137343f
C1564 uio_oe[5] VGND 0.137343f
C1565 uio_oe[6] VGND 0.137343f
C1566 uio_oe[7] VGND 0.289256f
C1567 uio_in[6] VGND 19.971539f
C1568 uio_in[5] VGND 15.647288f
C1569 ui_in[0] VGND 14.124138f
C1570 ui_in[1] VGND 12.519364f
C1571 uio_in[1] VGND 15.046968f
C1572 uio_in[2] VGND 15.199068f
C1573 ui_in[2] VGND 11.54435f
C1574 ui_in[3] VGND 12.04699f
C1575 uio_in[3] VGND 14.21004f
C1576 uio_in[4] VGND 14.381983f
C1577 uio_in[0] VGND 15.490564f
C1578 ui_in[7] VGND 15.539585f
C1579 ui_in[6] VGND 12.882964f
C1580 ui_in[5] VGND 10.864614f
C1581 ui_in[4] VGND 9.591749f
C1582 uo_out[0] VGND 9.065311f
C1583 uo_out[1] VGND 8.284716f
C1584 uo_out[2] VGND 7.409694f
C1585 uo_out[3] VGND 5.486512f
C1586 uo_out[4] VGND 3.7559f
C1587 uo_out[5] VGND 3.29391f
C1588 uo_out[6] VGND 2.83951f
C1589 uo_out[7] VGND 2.66217f
C1590 ua[0] VGND 9.46517f
C1591 VDPWR VGND 0.356001p
C1592 a_25284_5108# VGND 0.372398f
C1593 a_16786_5138# VGND 0.371932f
C1594 input_stage_andpwr_0.nand_gate_0.out VGND 0.873125f
C1595 input_stage_0.nand_gate_0.out VGND 0.872787f
C1596 a_24790_6672# VGND 0.387205f
C1597 a_24790_6936# VGND 0.612975f
C1598 input_stage_andpwr_0.fine_delay_unit_0.in VGND 1.81838f
C1599 a_23820_7082# VGND 0.731446f
C1600 a_16292_6702# VGND 0.387205f
C1601 a_16292_6966# VGND 0.612975f
C1602 input_stage_0.fine_delay_unit_0.in VGND 1.8013f
C1603 a_15322_7112# VGND 0.731446f
C1604 a_24790_8050# VGND 0.387205f
C1605 a_24790_8314# VGND 0.612975f
C1606 input_stage_andpwr_0.fine_delay_unit_1.in VGND 1.68519f
C1607 a_23820_8460# VGND 0.739963f
C1608 a_16292_8080# VGND 0.387205f
C1609 a_16292_8344# VGND 0.612975f
C1610 input_stage_0.fine_delay_unit_1.in VGND 1.67858f
C1611 a_15322_8490# VGND 0.739963f
C1612 variable_delay_short_0.in VGND 1.97381f
C1613 variable_delay_dummy_0.in VGND 1.96449f
C1614 a_25060_11366# VGND 0.71648f
C1615 a_24240_11366# VGND 0.037888f
C1616 a_16500_11634# VGND 0.71648f
C1617 a_15680_11634# VGND 0.037888f
C1618 a_7140_10670# VGND 1.49885f
C1619 a_25060_12248# VGND 0.717347f
C1620 a_24240_12248# VGND 0.043128f
C1621 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en VGND 2.516856f
C1622 variable_delay_dummy_0.out VGND 5.71113f
C1623 a_16500_12516# VGND 0.717347f
C1624 a_15680_12516# VGND 0.043128f
C1625 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en VGND 2.851508f
C1626 variable_delay_short_0.variable_delay_unit_1.in VGND 3.604031f
C1627 variable_delay_short_0.out VGND 8.859031f
C1628 variable_delay_dummy_0.variable_delay_unit_1.in VGND 4.168124f
C1629 a_9330_13764# VGND 0.629875f
C1630 a_25060_14314# VGND 0.71648f
C1631 a_24240_14314# VGND 0.037888f
C1632 a_9330_14054# VGND 0.622523f
C1633 tdc_0.start_buffer_0.start_delay VGND 3.694501f
C1634 tdc_0.start_buffer_0.start_buff VGND 5.257338f
C1635 a_16500_14582# VGND 0.71648f
C1636 a_15680_14582# VGND 0.037888f
C1637 variable_delay_dummy_0.variable_delay_unit_1.forward VGND 2.636476f
C1638 a_9330_14344# VGND 0.622523f
C1639 a_9330_14634# VGND 0.622248f
C1640 variable_delay_short_0.variable_delay_unit_1.out VGND 2.21957f
C1641 a_25060_15196# VGND 0.717347f
C1642 a_24240_15196# VGND 0.043128f
C1643 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en VGND 2.517556f
C1644 a_9330_14924# VGND 0.622523f
C1645 variable_delay_dummy_0.variable_delay_unit_1.out VGND 2.29732f
C1646 a_16500_15464# VGND 0.784074f
C1647 a_15680_15464# VGND 0.114203f
C1648 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en VGND 2.963248f
C1649 a_9330_15214# VGND 0.622289f
C1650 a_9330_15504# VGND 0.622536f
C1651 tdc_0.diff_gen_0.delay_unit_2_1.in_2 VGND 3.077349f
C1652 tdc_0.diff_gen_0.delay_unit_2_1.in_1 VGND 2.012721f
C1653 variable_delay_short_0.variable_delay_unit_2.in VGND 3.604041f
C1654 a_9330_15794# VGND 1.49187f
C1655 tdc_0.diff_gen_0.delay_unit_2_2.in_2 VGND 3.163373f
C1656 tdc_0.diff_gen_0.delay_unit_2_2.in_1 VGND 2.006561f
C1657 a_25060_17262# VGND 0.71648f
C1658 a_24240_17262# VGND 0.037888f
C1659 variable_delay_short_0.variable_delay_unit_2.out VGND 2.21957f
C1660 a_25060_18144# VGND 0.717347f
C1661 a_24240_18144# VGND 0.043128f
C1662 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en VGND 2.517556f
C1663 tdc_0.diff_gen_0.delay_unit_2_3.in_2 VGND 3.077369f
C1664 tdc_0.diff_gen_0.delay_unit_2_3.in_1 VGND 2.006501f
C1665 variable_delay_short_0.variable_delay_unit_3.in VGND 3.604041f
C1666 tdc_0.diff_gen_0.delay_unit_2_4.in_2 VGND 3.163433f
C1667 tdc_0.diff_gen_0.delay_unit_2_4.in_1 VGND 2.006681f
C1668 a_25060_20210# VGND 0.71648f
C1669 a_24240_20210# VGND 0.037888f
C1670 tdc_0.diff_gen_0.delay_unit_2_5.in_2 VGND 3.163143f
C1671 variable_delay_short_0.variable_delay_unit_3.out VGND 2.21957f
C1672 a_25060_21092# VGND 0.717347f
C1673 a_24240_21092# VGND 0.043128f
C1674 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en VGND 2.517556f
C1675 tdc_0.diff_gen_0.delay_unit_2_6.in_2 VGND 3.083859f
C1676 tdc_0.diff_gen_0.delay_unit_2_6.in_1 VGND 2.070971f
C1677 variable_delay_short_0.variable_delay_unit_4.in VGND 3.604041f
C1678 a_25060_23158# VGND 0.71648f
C1679 a_24240_23158# VGND 0.037888f
C1680 variable_delay_short_0.variable_delay_unit_4.out VGND 2.21957f
C1681 a_25060_24040# VGND 0.717347f
C1682 a_24240_24040# VGND 0.043128f
C1683 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en VGND 2.517556f
C1684 a_13254_23752# VGND 0.190873f
C1685 a_12310_23706# VGND 0.838649f
C1686 a_12420_23752# VGND 0.024712f
C1687 a_13254_24130# VGND 0.192269f
C1688 a_12420_24130# VGND 0.023462f
C1689 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VGND 0.583709f
C1690 a_12308_24168# VGND 0.823328f
C1691 a_10108_23452# VGND 0.354057f
C1692 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VGND 6.034074f
C1693 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VGND 7.095738f
C1694 tdc_0.vernier_delay_line_0.start_neg VGND 3.594784f
C1695 tdc_0.vernier_delay_line_0.start_pos VGND 2.750328f
C1696 variable_delay_short_0.variable_delay_unit_5.in VGND 3.860429f
C1697 a_25060_26106# VGND 0.71648f
C1698 a_24240_26106# VGND 0.037888f
C1699 variable_delay_short_0.variable_delay_unit_5.forward VGND 2.636476f
C1700 a_13254_26034# VGND 0.190624f
C1701 a_12310_25988# VGND 0.829382f
C1702 a_12420_26034# VGND 0.024712f
C1703 a_13254_26412# VGND 0.192129f
C1704 a_12420_26412# VGND 0.023462f
C1705 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VGND 0.583105f
C1706 a_12308_26450# VGND 0.823144f
C1707 variable_delay_short_0.variable_delay_unit_5.out VGND 2.29732f
C1708 a_25060_26988# VGND 0.784074f
C1709 a_24240_26988# VGND 0.114203f
C1710 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en VGND 2.963248f
C1711 a_10108_25734# VGND 0.354057f
C1712 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1713 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1714 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 VGND 6.192364f
C1715 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 VGND 5.851951f
C1716 a_13254_28316# VGND 0.190624f
C1717 a_12310_28270# VGND 0.829382f
C1718 a_12420_28316# VGND 0.024712f
C1719 a_13254_28694# VGND 0.192129f
C1720 a_12420_28694# VGND 0.023462f
C1721 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VGND 0.583105f
C1722 a_12308_28732# VGND 0.823144f
C1723 a_10108_28016# VGND 0.354057f
C1724 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1725 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1726 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 VGND 6.192265f
C1727 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 VGND 5.68077f
C1728 a_13254_30598# VGND 0.190624f
C1729 a_12310_30552# VGND 0.829382f
C1730 a_12420_30598# VGND 0.024712f
C1731 a_13254_30976# VGND 0.192129f
C1732 a_12420_30976# VGND 0.023462f
C1733 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VGND 0.583105f
C1734 a_12308_31014# VGND 0.823144f
C1735 a_10108_30298# VGND 0.354057f
C1736 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1737 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1738 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VGND 6.192265f
C1739 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VGND 5.68077f
C1740 a_13254_32880# VGND 0.190624f
C1741 a_12310_32834# VGND 0.829382f
C1742 a_12420_32880# VGND 0.024712f
C1743 a_13254_33258# VGND 0.192129f
C1744 a_12420_33258# VGND 0.023462f
C1745 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VGND 0.583105f
C1746 a_12308_33296# VGND 0.823144f
C1747 a_10108_32580# VGND 0.354057f
C1748 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1749 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1750 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 VGND 6.021708f
C1751 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 VGND 5.489025f
C1752 a_13254_35162# VGND 0.190624f
C1753 a_12310_35116# VGND 0.829382f
C1754 a_12420_35162# VGND 0.024712f
C1755 a_13254_35540# VGND 0.192129f
C1756 a_12420_35540# VGND 0.023462f
C1757 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VGND 0.583105f
C1758 a_12308_35578# VGND 0.823144f
C1759 a_10108_34862# VGND 0.354057f
C1760 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1761 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1762 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 VGND 6.021708f
C1763 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 VGND 5.489025f
C1764 a_13254_37444# VGND 0.190624f
C1765 a_12310_37398# VGND 0.829382f
C1766 a_12420_37444# VGND 0.024712f
C1767 a_13254_37822# VGND 0.192129f
C1768 a_12420_37822# VGND 0.023462f
C1769 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VGND 0.583105f
C1770 a_12308_37860# VGND 0.823144f
C1771 a_10108_37144# VGND 0.354057f
C1772 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1773 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1774 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 VGND 6.192265f
C1775 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 VGND 5.68077f
C1776 a_13254_39726# VGND 0.190624f
C1777 a_12310_39680# VGND 0.829382f
C1778 a_12420_39726# VGND 0.024712f
C1779 a_13254_40104# VGND 0.192129f
C1780 a_12420_40104# VGND 0.023462f
C1781 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VGND 0.583308f
C1782 a_12308_40142# VGND 0.830326f
C1783 a_10108_39426# VGND 0.354057f
C1784 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VGND 6.505114f
C1785 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VGND 6.446748f
C1786 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 VGND 6.192265f
C1787 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 VGND 5.68077f
C1788 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 VGND 0.974288f
C1789 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VGND 1.24637f
C1790 uio_in[2].t0 VGND 0.083134f
C1791 uio_in[2].n0 VGND 7.1868f
C1792 ui_in[1].t0 VGND 0.062351f
C1793 ui_in[1].n0 VGND 4.87703f
C1794 uio_in[5].t0 VGND 0.045056f
C1795 uio_in[5].t1 VGND 0.06074f
C1796 uio_in[5].n0 VGND 0.067592f
C1797 uio_in[5].n1 VGND 4.90746f
C1798 uio_in[4].t0 VGND 0.084602f
C1799 uio_in[4].n0 VGND 6.89354f
C1800 uio_in[1].t0 VGND 0.064466f
C1801 uio_in[1].n0 VGND 6.45166f
C1802 ui_in[3].t0 VGND 0.046163f
C1803 ui_in[3].n0 VGND 3.40417f
C1804 variable_delay_short_0.variable_delay_unit_1.in.t4 VGND 0.017058f
C1805 variable_delay_short_0.variable_delay_unit_1.in.t5 VGND 0.044984f
C1806 variable_delay_short_0.variable_delay_unit_1.in.n0 VGND 0.04731f
C1807 variable_delay_short_0.variable_delay_unit_1.in.t0 VGND 0.033139f
C1808 variable_delay_short_0.variable_delay_unit_1.in.t1 VGND 0.105354f
C1809 variable_delay_short_0.variable_delay_unit_1.in.n1 VGND 0.255341f
C1810 variable_delay_short_0.variable_delay_unit_1.in.t2 VGND 0.042943f
C1811 variable_delay_short_0.variable_delay_unit_1.in.t3 VGND 0.013862f
C1812 variable_delay_short_0.variable_delay_unit_1.in.n2 VGND 0.045161f
C1813 variable_delay_short_0.variable_delay_unit_1.in.n3 VGND 0.418008f
C1814 variable_delay_short_0.variable_delay_unit_2.in.t4 VGND 0.017058f
C1815 variable_delay_short_0.variable_delay_unit_2.in.t5 VGND 0.044984f
C1816 variable_delay_short_0.variable_delay_unit_2.in.n0 VGND 0.04731f
C1817 variable_delay_short_0.variable_delay_unit_2.in.t1 VGND 0.033139f
C1818 variable_delay_short_0.variable_delay_unit_2.in.t0 VGND 0.105354f
C1819 variable_delay_short_0.variable_delay_unit_2.in.n1 VGND 0.255341f
C1820 variable_delay_short_0.variable_delay_unit_2.in.t2 VGND 0.042943f
C1821 variable_delay_short_0.variable_delay_unit_2.in.t3 VGND 0.013862f
C1822 variable_delay_short_0.variable_delay_unit_2.in.n2 VGND 0.045161f
C1823 variable_delay_short_0.variable_delay_unit_2.in.n3 VGND 0.418008f
C1824 a_10108_37672.t3 VGND 0.059028f
C1825 a_10108_37672.t2 VGND 0.059028f
C1826 a_10108_37672.t5 VGND 0.059028f
C1827 a_10108_37672.n0 VGND 0.136068f
C1828 a_10108_37672.t0 VGND 0.059028f
C1829 a_10108_37672.t1 VGND 0.059028f
C1830 a_10108_37672.n1 VGND 0.139449f
C1831 a_10108_37672.n2 VGND 1.11221f
C1832 a_10108_37672.n3 VGND 0.258102f
C1833 a_10108_37672.t4 VGND 0.059028f
C1834 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 VGND 0.930597f
C1835 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.765644f
C1836 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.087567f
C1837 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C1838 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C1839 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C1840 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C1841 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C1842 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C1843 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.089004f
C1844 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C1845 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C1846 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C1847 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C1848 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C1849 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C1850 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C1851 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 VGND 0.748416f
C1852 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C1853 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C1854 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.096169f
C1855 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C1856 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C1857 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C1858 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C1859 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C1860 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C1861 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C1862 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C1863 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C1864 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C1865 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C1866 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C1867 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C1868 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C1869 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C1870 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C1871 ui_in[0].t0 VGND 0.028496f
C1872 ui_in[0].n0 VGND 2.53887f
C1873 uio_in[3].t0 VGND 0.07563f
C1874 uio_in[3].n0 VGND 7.04584f
C1875 uo_out[2].t5 VGND 0.01472f
C1876 uo_out[2].t4 VGND 0.04976f
C1877 uo_out[2].n0 VGND 0.040339f
C1878 uo_out[2].t3 VGND 0.028671f
C1879 uo_out[2].t1 VGND 0.028671f
C1880 uo_out[2].n1 VGND 0.060931f
C1881 uo_out[2].n2 VGND 0.265829f
C1882 uo_out[2].t0 VGND 0.009557f
C1883 uo_out[2].t2 VGND 0.009557f
C1884 uo_out[2].n3 VGND 0.020748f
C1885 uo_out[2].n4 VGND 0.070592f
C1886 uo_out[2].n5 VGND 1.57081f
C1887 uo_out[1].t5 VGND 0.015076f
C1888 uo_out[1].t4 VGND 0.050965f
C1889 uo_out[1].n0 VGND 0.041315f
C1890 uo_out[1].t1 VGND 0.029365f
C1891 uo_out[1].t3 VGND 0.029365f
C1892 uo_out[1].n1 VGND 0.062406f
C1893 uo_out[1].n2 VGND 0.272264f
C1894 uo_out[1].t2 VGND 0.009788f
C1895 uo_out[1].t0 VGND 0.009788f
C1896 uo_out[1].n3 VGND 0.02125f
C1897 uo_out[1].n4 VGND 0.072301f
C1898 uo_out[1].n5 VGND 1.84327f
C1899 ui_in[2].t0 VGND 0.055937f
C1900 ui_in[2].n0 VGND 4.70026f
C1901 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 VGND 0.020532f
C1902 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 VGND 0.020532f
C1903 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 VGND 0.048092f
C1904 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 VGND 0.061597f
C1905 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 VGND 0.061597f
C1906 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 VGND 0.125485f
C1907 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 VGND 0.522094f
C1908 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 VGND 0.075157f
C1909 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 VGND 0.227425f
C1910 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 VGND 0.55466f
C1911 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 VGND 0.283681f
C1912 variable_delay_dummy_0.variable_delay_unit_1.forward.t3 VGND 0.025654f
C1913 variable_delay_dummy_0.variable_delay_unit_1.forward.t2 VGND 0.067654f
C1914 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 VGND 0.071153f
C1915 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 VGND 0.04984f
C1916 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 VGND 0.15845f
C1917 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 VGND 0.384027f
C1918 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 VGND 0.628675f
C1919 variable_delay_dummy_0.variable_delay_unit_1.in.t5 VGND 0.025993f
C1920 variable_delay_dummy_0.variable_delay_unit_1.in.t4 VGND 0.068546f
C1921 variable_delay_dummy_0.variable_delay_unit_1.in.n0 VGND 0.072091f
C1922 variable_delay_dummy_0.variable_delay_unit_1.in.t0 VGND 0.050497f
C1923 variable_delay_dummy_0.variable_delay_unit_1.in.t1 VGND 0.160539f
C1924 variable_delay_dummy_0.variable_delay_unit_1.in.n1 VGND 0.389091f
C1925 variable_delay_dummy_0.variable_delay_unit_1.in.t3 VGND 0.065437f
C1926 variable_delay_dummy_0.variable_delay_unit_1.in.t2 VGND 0.021123f
C1927 variable_delay_dummy_0.variable_delay_unit_1.in.n2 VGND 0.068816f
C1928 variable_delay_dummy_0.variable_delay_unit_1.in.n3 VGND 0.636965f
C1929 a_10108_33108.t2 VGND 0.059028f
C1930 a_10108_33108.t1 VGND 0.059028f
C1931 a_10108_33108.t0 VGND 0.059028f
C1932 a_10108_33108.n0 VGND 0.139449f
C1933 a_10108_33108.t3 VGND 0.059028f
C1934 a_10108_33108.t5 VGND 0.059028f
C1935 a_10108_33108.n1 VGND 0.258102f
C1936 a_10108_33108.n2 VGND 1.11221f
C1937 a_10108_33108.n3 VGND 0.136068f
C1938 a_10108_33108.t4 VGND 0.059028f
C1939 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 VGND 0.09757f
C1940 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 VGND 0.030153f
C1941 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 VGND 0.265657f
C1942 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 VGND 0.039259f
C1943 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 VGND 0.012524f
C1944 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 VGND 0.027534f
C1945 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 VGND 0.039259f
C1946 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 VGND 0.012524f
C1947 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 VGND 0.027357f
C1948 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 VGND 0.008823f
C1949 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VGND 0.039259f
C1950 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 VGND 0.012524f
C1951 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 VGND 0.027534f
C1952 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 VGND 0.039259f
C1953 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 VGND 0.012524f
C1954 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 VGND 0.027357f
C1955 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 VGND 0.008728f
C1956 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 VGND 0.135162f
C1957 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 VGND 0.046129f
C1958 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 VGND 0.046129f
C1959 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 VGND 0.054044f
C1960 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 VGND 0.046129f
C1961 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 VGND 0.046129f
C1962 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 VGND 0.0538f
C1963 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 VGND 0.495704f
C1964 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 VGND 0.119944f
C1965 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 VGND 0.025758f
C1966 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 VGND 0.025758f
C1967 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 VGND 0.055083f
C1968 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VGND 0.008586f
C1969 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 VGND 0.008586f
C1970 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 VGND 0.01864f
C1971 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 VGND 0.221512f
C1972 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 VGND 0.09757f
C1973 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 VGND 0.030153f
C1974 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 VGND 0.234486f
C1975 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 VGND 0.050613f
C1976 tdc_0.vernier_delay_line_0.start_neg.t1 VGND 0.153672f
C1977 tdc_0.vernier_delay_line_0.start_neg.t0 VGND 0.047491f
C1978 tdc_0.vernier_delay_line_0.start_neg.n0 VGND 0.42006f
C1979 tdc_0.vernier_delay_line_0.start_neg.t8 VGND 0.061832f
C1980 tdc_0.vernier_delay_line_0.start_neg.t15 VGND 0.019725f
C1981 tdc_0.vernier_delay_line_0.start_neg.n1 VGND 0.043367f
C1982 tdc_0.vernier_delay_line_0.start_neg.t14 VGND 0.061832f
C1983 tdc_0.vernier_delay_line_0.start_neg.t13 VGND 0.019725f
C1984 tdc_0.vernier_delay_line_0.start_neg.n2 VGND 0.043087f
C1985 tdc_0.vernier_delay_line_0.start_neg.n3 VGND 0.013896f
C1986 tdc_0.vernier_delay_line_0.start_neg.t12 VGND 0.061832f
C1987 tdc_0.vernier_delay_line_0.start_neg.t10 VGND 0.019725f
C1988 tdc_0.vernier_delay_line_0.start_neg.n4 VGND 0.043367f
C1989 tdc_0.vernier_delay_line_0.start_neg.t11 VGND 0.061832f
C1990 tdc_0.vernier_delay_line_0.start_neg.t9 VGND 0.019725f
C1991 tdc_0.vernier_delay_line_0.start_neg.n5 VGND 0.043087f
C1992 tdc_0.vernier_delay_line_0.start_neg.n6 VGND 0.013747f
C1993 tdc_0.vernier_delay_line_0.start_neg.n7 VGND 0.187263f
C1994 tdc_0.vernier_delay_line_0.start_neg.t5 VGND 0.040569f
C1995 tdc_0.vernier_delay_line_0.start_neg.t6 VGND 0.040569f
C1996 tdc_0.vernier_delay_line_0.start_neg.n8 VGND 0.086755f
C1997 tdc_0.vernier_delay_line_0.start_neg.t3 VGND 0.013523f
C1998 tdc_0.vernier_delay_line_0.start_neg.t4 VGND 0.013523f
C1999 tdc_0.vernier_delay_line_0.start_neg.n9 VGND 0.029358f
C2000 tdc_0.vernier_delay_line_0.start_neg.n10 VGND 0.348878f
C2001 tdc_0.vernier_delay_line_0.start_neg.t7 VGND 0.153672f
C2002 tdc_0.vernier_delay_line_0.start_neg.t2 VGND 0.047491f
C2003 tdc_0.vernier_delay_line_0.start_neg.n11 VGND 0.369312f
C2004 tdc_0.vernier_delay_line_0.start_neg.n12 VGND 0.079715f
C2005 uio_in[0].t1 VGND 0.072685f
C2006 uio_in[0].t5 VGND 0.078634f
C2007 uio_in[0].n0 VGND 0.077149f
C2008 uio_in[0].t7 VGND 0.078369f
C2009 uio_in[0].n1 VGND 0.053689f
C2010 uio_in[0].t0 VGND 0.022787f
C2011 uio_in[0].t2 VGND 0.029248f
C2012 uio_in[0].t6 VGND 0.029248f
C2013 uio_in[0].n2 VGND 0.087662f
C2014 uio_in[0].n3 VGND 0.531341f
C2015 uio_in[0].n4 VGND 5.469f
C2016 uio_in[0].t3 VGND 0.073684f
C2017 uio_in[0].t4 VGND 0.023785f
C2018 uio_in[0].n5 VGND 0.074548f
C2019 uio_in[0].n6 VGND 0.62346f
C2020 uio_in[6].t0 VGND 0.019238f
C2021 uio_in[6].t2 VGND 0.028339f
C2022 uio_in[6].n0 VGND 0.0304f
C2023 uio_in[6].t1 VGND 0.019238f
C2024 uio_in[6].t3 VGND 0.028339f
C2025 uio_in[6].n1 VGND 0.0304f
C2026 uio_in[6].n2 VGND 3.91151f
C2027 ui_in[6].t0 VGND 0.064986f
C2028 ui_in[6].t1 VGND 0.070305f
C2029 ui_in[6].n0 VGND 0.068977f
C2030 ui_in[6].t5 VGND 0.070068f
C2031 ui_in[6].n1 VGND 0.048001f
C2032 ui_in[6].t6 VGND 0.020373f
C2033 ui_in[6].t7 VGND 0.02615f
C2034 ui_in[6].t4 VGND 0.02615f
C2035 ui_in[6].n2 VGND 0.078377f
C2036 ui_in[6].n3 VGND 0.397332f
C2037 ui_in[6].n4 VGND 4.07223f
C2038 ui_in[6].t2 VGND 0.065879f
C2039 ui_in[6].t3 VGND 0.021265f
C2040 ui_in[6].n5 VGND 0.066651f
C2041 ui_in[6].n6 VGND 0.565747f
C2042 ui_in[7].t1 VGND 0.08368f
C2043 ui_in[7].t5 VGND 0.090529f
C2044 ui_in[7].n0 VGND 0.088818f
C2045 ui_in[7].t7 VGND 0.090223f
C2046 ui_in[7].n1 VGND 0.06181f
C2047 ui_in[7].t0 VGND 0.026234f
C2048 ui_in[7].t4 VGND 0.033672f
C2049 ui_in[7].t6 VGND 0.033672f
C2050 ui_in[7].n2 VGND 0.100922f
C2051 ui_in[7].n3 VGND 0.609031f
C2052 ui_in[7].n4 VGND 5.81591f
C2053 ui_in[7].t2 VGND 0.084829f
C2054 ui_in[7].t3 VGND 0.027383f
C2055 ui_in[7].n5 VGND 0.085824f
C2056 ui_in[7].n6 VGND 0.719999f
C2057 tdc_0.vernier_delay_line_0.start_pos.t11 VGND 0.086445f
C2058 tdc_0.vernier_delay_line_0.start_pos.t9 VGND 0.027576f
C2059 tdc_0.vernier_delay_line_0.start_pos.n0 VGND 0.060238f
C2060 tdc_0.vernier_delay_line_0.start_pos.t8 VGND 0.086445f
C2061 tdc_0.vernier_delay_line_0.start_pos.t15 VGND 0.027576f
C2062 tdc_0.vernier_delay_line_0.start_pos.n1 VGND 0.060629f
C2063 tdc_0.vernier_delay_line_0.start_pos.n2 VGND 0.01943f
C2064 tdc_0.vernier_delay_line_0.start_pos.t14 VGND 0.086445f
C2065 tdc_0.vernier_delay_line_0.start_pos.t13 VGND 0.027576f
C2066 tdc_0.vernier_delay_line_0.start_pos.n3 VGND 0.060629f
C2067 tdc_0.vernier_delay_line_0.start_pos.t12 VGND 0.086445f
C2068 tdc_0.vernier_delay_line_0.start_pos.t10 VGND 0.027576f
C2069 tdc_0.vernier_delay_line_0.start_pos.n4 VGND 0.060238f
C2070 tdc_0.vernier_delay_line_0.start_pos.n5 VGND 0.019219f
C2071 tdc_0.vernier_delay_line_0.start_pos.n6 VGND 0.507295f
C2072 tdc_0.vernier_delay_line_0.start_pos.t6 VGND 0.069183f
C2073 tdc_0.vernier_delay_line_0.start_pos.t7 VGND 0.209408f
C2074 tdc_0.vernier_delay_line_0.start_pos.n7 VGND 0.531486f
C2075 tdc_0.vernier_delay_line_0.start_pos.n8 VGND 0.276923f
C2076 tdc_0.vernier_delay_line_0.start_pos.t1 VGND 0.018906f
C2077 tdc_0.vernier_delay_line_0.start_pos.t2 VGND 0.018906f
C2078 tdc_0.vernier_delay_line_0.start_pos.n9 VGND 0.044282f
C2079 tdc_0.vernier_delay_line_0.start_pos.t3 VGND 0.056718f
C2080 tdc_0.vernier_delay_line_0.start_pos.t4 VGND 0.056718f
C2081 tdc_0.vernier_delay_line_0.start_pos.n10 VGND 0.115544f
C2082 tdc_0.vernier_delay_line_0.start_pos.n11 VGND 0.480734f
C2083 tdc_0.vernier_delay_line_0.start_pos.t0 VGND 0.069203f
C2084 tdc_0.vernier_delay_line_0.start_pos.t5 VGND 0.209408f
C2085 tdc_0.vernier_delay_line_0.start_pos.n12 VGND 0.51072f
C2086 tdc_0.vernier_delay_line_0.start_pos.n13 VGND 0.261208f
C2087 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 VGND 0.165681f
C2088 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 VGND 0.051203f
C2089 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 VGND 0.451103f
C2090 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 VGND 0.066664f
C2091 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 VGND 0.021266f
C2092 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 VGND 0.046756f
C2093 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 VGND 0.066664f
C2094 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 VGND 0.021266f
C2095 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 VGND 0.046454f
C2096 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 VGND 0.014982f
C2097 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 VGND 0.066664f
C2098 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 VGND 0.021266f
C2099 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 VGND 0.046756f
C2100 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 VGND 0.066664f
C2101 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 VGND 0.021266f
C2102 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 VGND 0.046454f
C2103 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 VGND 0.014821f
C2104 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 VGND 0.229513f
C2105 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 VGND 0.043739f
C2106 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 VGND 0.043739f
C2107 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 VGND 0.093535f
C2108 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 VGND 0.01458f
C2109 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 VGND 0.01458f
C2110 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 VGND 0.031652f
C2111 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 VGND 0.376142f
C2112 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 VGND 0.165681f
C2113 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 VGND 0.051203f
C2114 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 VGND 0.398173f
C2115 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 VGND 0.085944f
C2116 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VGND 0.059856f
C2117 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 VGND 0.019094f
C2118 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2119 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2120 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 VGND 0.019094f
C2121 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2122 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2123 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 VGND 0.059856f
C2124 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VGND 0.019094f
C2125 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2126 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 VGND 0.059856f
C2127 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 VGND 0.019094f
C2128 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2129 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2130 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2131 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VGND 0.047903f
C2132 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VGND 0.144997f
C2133 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2134 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 VGND 0.191745f
C2135 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VGND 0.013091f
C2136 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 VGND 0.013091f
C2137 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 VGND 0.030662f
C2138 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 VGND 0.039272f
C2139 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 VGND 0.039272f
C2140 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 VGND 0.080004f
C2141 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 VGND 0.332866f
C2142 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 VGND 0.060722f
C2143 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2144 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 VGND 0.070899f
C2145 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 VGND 0.060722f
C2146 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 VGND 0.060722f
C2147 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 VGND 0.070523f
C2148 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 VGND 0.632153f
C2149 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 VGND 0.045973f
C2150 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 VGND 0.156775f
C2151 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 VGND 0.144997f
C2152 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 VGND 0.240639f
C2153 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 VGND 0.180864f
C2154 ui_in[4].t3 VGND 0.039584f
C2155 ui_in[4].t5 VGND 0.012778f
C2156 ui_in[4].n0 VGND 0.040049f
C2157 ui_in[4].t0 VGND 0.039048f
C2158 ui_in[4].t2 VGND 0.042244f
C2159 ui_in[4].n1 VGND 0.041446f
C2160 ui_in[4].t6 VGND 0.042102f
C2161 ui_in[4].n2 VGND 0.028843f
C2162 ui_in[4].t7 VGND 0.012242f
C2163 ui_in[4].t1 VGND 0.015712f
C2164 ui_in[4].t4 VGND 0.015712f
C2165 ui_in[4].n3 VGND 0.047094f
C2166 ui_in[4].n4 VGND 0.28086f
C2167 ui_in[4].n5 VGND 1.95509f
C2168 ui_in[4].n6 VGND 0.343484f
C2169 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 VGND 0.059856f
C2170 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 VGND 0.019094f
C2171 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2172 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 VGND 0.059856f
C2173 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2174 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2175 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2176 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 VGND 0.059856f
C2177 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 VGND 0.019094f
C2178 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2179 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2180 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2181 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2182 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2183 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2184 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 VGND 0.047903f
C2185 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 VGND 0.144997f
C2186 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2187 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 VGND 0.013091f
C2188 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 VGND 0.013091f
C2189 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 VGND 0.030662f
C2190 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VGND 0.039272f
C2191 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 VGND 0.039272f
C2192 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 VGND 0.080004f
C2193 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 VGND 0.332866f
C2194 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 VGND 0.060722f
C2195 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 VGND 0.060722f
C2196 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 VGND 0.070899f
C2197 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2198 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 VGND 0.060722f
C2199 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 VGND 0.070523f
C2200 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 VGND 0.632153f
C2201 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 VGND 0.045973f
C2202 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 VGND 0.156775f
C2203 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 VGND 0.144997f
C2204 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 VGND 0.240639f
C2205 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 VGND 0.180864f
C2206 variable_delay_short_0.variable_delay_unit_4.in.t4 VGND 0.017058f
C2207 variable_delay_short_0.variable_delay_unit_4.in.t5 VGND 0.044984f
C2208 variable_delay_short_0.variable_delay_unit_4.in.n0 VGND 0.04731f
C2209 variable_delay_short_0.variable_delay_unit_4.in.t0 VGND 0.033139f
C2210 variable_delay_short_0.variable_delay_unit_4.in.t1 VGND 0.105354f
C2211 variable_delay_short_0.variable_delay_unit_4.in.n1 VGND 0.255341f
C2212 variable_delay_short_0.variable_delay_unit_4.in.t2 VGND 0.042943f
C2213 variable_delay_short_0.variable_delay_unit_4.in.t3 VGND 0.013862f
C2214 variable_delay_short_0.variable_delay_unit_4.in.n2 VGND 0.045161f
C2215 variable_delay_short_0.variable_delay_unit_4.in.n3 VGND 0.418008f
C2216 variable_delay_short_0.variable_delay_unit_3.in.t4 VGND 0.017058f
C2217 variable_delay_short_0.variable_delay_unit_3.in.t5 VGND 0.044984f
C2218 variable_delay_short_0.variable_delay_unit_3.in.n0 VGND 0.04731f
C2219 variable_delay_short_0.variable_delay_unit_3.in.t0 VGND 0.033139f
C2220 variable_delay_short_0.variable_delay_unit_3.in.t1 VGND 0.105354f
C2221 variable_delay_short_0.variable_delay_unit_3.in.n1 VGND 0.255341f
C2222 variable_delay_short_0.variable_delay_unit_3.in.t2 VGND 0.042943f
C2223 variable_delay_short_0.variable_delay_unit_3.in.t3 VGND 0.013862f
C2224 variable_delay_short_0.variable_delay_unit_3.in.n2 VGND 0.045161f
C2225 variable_delay_short_0.variable_delay_unit_3.in.n3 VGND 0.418008f
C2226 a_10108_23980.t2 VGND 0.059028f
C2227 a_10108_23980.t0 VGND 0.059028f
C2228 a_10108_23980.t1 VGND 0.059028f
C2229 a_10108_23980.n0 VGND 0.139449f
C2230 a_10108_23980.t3 VGND 0.059028f
C2231 a_10108_23980.t5 VGND 0.059028f
C2232 a_10108_23980.n1 VGND 0.258102f
C2233 a_10108_23980.n2 VGND 1.11221f
C2234 a_10108_23980.n3 VGND 0.136068f
C2235 a_10108_23980.t4 VGND 0.059028f
C2236 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 VGND 0.09757f
C2237 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 VGND 0.030153f
C2238 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2239 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VGND 0.039259f
C2240 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2241 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2242 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 VGND 0.039259f
C2243 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 VGND 0.012524f
C2244 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2245 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2246 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 VGND 0.039259f
C2247 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2248 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2249 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2250 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 VGND 0.012524f
C2251 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2252 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2253 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2254 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 VGND 0.046129f
C2255 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 VGND 0.046129f
C2256 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2257 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 VGND 0.046129f
C2258 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 VGND 0.046129f
C2259 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2260 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2261 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 VGND 0.025758f
C2262 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 VGND 0.025758f
C2263 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2264 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VGND 0.008586f
C2265 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 VGND 0.008586f
C2266 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2267 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2268 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 VGND 0.09757f
C2269 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 VGND 0.030153f
C2270 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2271 a_10958_30210.t3 VGND 0.024913f
C2272 a_10958_30210.t0 VGND 0.024913f
C2273 a_10958_30210.t2 VGND 0.024913f
C2274 a_10958_30210.n0 VGND 0.059872f
C2275 a_10958_30210.t12 VGND 0.096748f
C2276 a_10958_30210.t5 VGND 0.024913f
C2277 a_10958_30210.t9 VGND 0.024913f
C2278 a_10958_30210.n1 VGND 0.060504f
C2279 a_10958_30210.n2 VGND 0.369187f
C2280 a_10958_30210.t11 VGND 0.024913f
C2281 a_10958_30210.t7 VGND 0.024913f
C2282 a_10958_30210.n3 VGND 0.060504f
C2283 a_10958_30210.n4 VGND 0.182084f
C2284 a_10958_30210.t8 VGND 0.024913f
C2285 a_10958_30210.t10 VGND 0.024913f
C2286 a_10958_30210.n5 VGND 0.060504f
C2287 a_10958_30210.n6 VGND 0.221492f
C2288 a_10958_30210.t1 VGND 0.024913f
C2289 a_10958_30210.t6 VGND 0.024913f
C2290 a_10958_30210.n7 VGND 0.052659f
C2291 a_10958_30210.n8 VGND 0.137512f
C2292 a_10958_30210.n9 VGND 0.342225f
C2293 a_10958_30210.n10 VGND 0.057757f
C2294 a_10958_30210.t4 VGND 0.024913f
C2295 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 VGND 0.059856f
C2296 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2297 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2298 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 VGND 0.059856f
C2299 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 VGND 0.019094f
C2300 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2301 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2302 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2303 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2304 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2305 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 VGND 0.059856f
C2306 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 VGND 0.019094f
C2307 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2308 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2309 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2310 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VGND 0.047903f
C2311 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VGND 0.144997f
C2312 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2313 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 VGND 0.013091f
C2314 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 VGND 0.013091f
C2315 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 VGND 0.030662f
C2316 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 VGND 0.039272f
C2317 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 VGND 0.039272f
C2318 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 VGND 0.080004f
C2319 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 VGND 0.332866f
C2320 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 VGND 0.060722f
C2321 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 VGND 0.060722f
C2322 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 VGND 0.070899f
C2323 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 VGND 0.060722f
C2324 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 VGND 0.060722f
C2325 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 VGND 0.070523f
C2326 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 VGND 0.632153f
C2327 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 VGND 0.045973f
C2328 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 VGND 0.156775f
C2329 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 VGND 0.144997f
C2330 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 VGND 0.240639f
C2331 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 VGND 0.180864f
C2332 variable_delay_short_0.variable_delay_unit_5.forward.t2 VGND 0.025654f
C2333 variable_delay_short_0.variable_delay_unit_5.forward.t3 VGND 0.067654f
C2334 variable_delay_short_0.variable_delay_unit_5.forward.n0 VGND 0.071153f
C2335 variable_delay_short_0.variable_delay_unit_5.forward.t0 VGND 0.04984f
C2336 variable_delay_short_0.variable_delay_unit_5.forward.t1 VGND 0.15845f
C2337 variable_delay_short_0.variable_delay_unit_5.forward.n1 VGND 0.384027f
C2338 variable_delay_short_0.variable_delay_unit_5.forward.n2 VGND 0.628675f
C2339 variable_delay_short_0.variable_delay_unit_5.in.t4 VGND 0.021119f
C2340 variable_delay_short_0.variable_delay_unit_5.in.t5 VGND 0.055694f
C2341 variable_delay_short_0.variable_delay_unit_5.in.n0 VGND 0.058574f
C2342 variable_delay_short_0.variable_delay_unit_5.in.t0 VGND 0.041029f
C2343 variable_delay_short_0.variable_delay_unit_5.in.t1 VGND 0.130438f
C2344 variable_delay_short_0.variable_delay_unit_5.in.n1 VGND 0.316137f
C2345 variable_delay_short_0.variable_delay_unit_5.in.t2 VGND 0.053167f
C2346 variable_delay_short_0.variable_delay_unit_5.in.t3 VGND 0.017162f
C2347 variable_delay_short_0.variable_delay_unit_5.in.n2 VGND 0.055913f
C2348 variable_delay_short_0.variable_delay_unit_5.in.n3 VGND 0.517534f
C2349 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C2350 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C2351 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.087567f
C2352 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.039734f
C2353 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C2354 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.089004f
C2355 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C2356 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C2357 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C2358 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C2359 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C2360 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C2361 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C2362 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C2363 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C2364 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C2365 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C2366 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 VGND 0.025758f
C2367 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 VGND 0.025758f
C2368 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 VGND 0.055083f
C2369 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2370 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 VGND 0.008586f
C2371 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 VGND 0.01864f
C2372 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 VGND 0.221512f
C2373 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 VGND 0.09757f
C2374 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 VGND 0.030153f
C2375 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 VGND 0.234486f
C2376 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 VGND 0.046129f
C2377 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2378 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 VGND 0.054044f
C2379 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 VGND 0.046129f
C2380 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2381 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 VGND 0.0538f
C2382 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 VGND 0.495704f
C2383 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 VGND 0.09757f
C2384 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 VGND 0.030153f
C2385 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 VGND 0.265657f
C2386 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VGND 0.039259f
C2387 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 VGND 0.012524f
C2388 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 VGND 0.027534f
C2389 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 VGND 0.039259f
C2390 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2391 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 VGND 0.027357f
C2392 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 VGND 0.008823f
C2393 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2394 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2395 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 VGND 0.027534f
C2396 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2397 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 VGND 0.012524f
C2398 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 VGND 0.027357f
C2399 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 VGND 0.008728f
C2400 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 VGND 0.135162f
C2401 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 VGND 0.086195f
C2402 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 VGND 0.027496f
C2403 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 VGND 0.060063f
C2404 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 VGND 0.086195f
C2405 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 VGND 0.027496f
C2406 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 VGND 0.060453f
C2407 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 VGND 0.019374f
C2408 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 VGND 0.086195f
C2409 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 VGND 0.027496f
C2410 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 VGND 0.060453f
C2411 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 VGND 0.086195f
C2412 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 VGND 0.027496f
C2413 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 VGND 0.060063f
C2414 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 VGND 0.019163f
C2415 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 VGND 0.505822f
C2416 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 VGND 0.068982f
C2417 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 VGND 0.2088f
C2418 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 VGND 0.529943f
C2419 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 VGND 0.27612f
C2420 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 VGND 0.018851f
C2421 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 VGND 0.018851f
C2422 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 VGND 0.044154f
C2423 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 VGND 0.056553f
C2424 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 VGND 0.056553f
C2425 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 VGND 0.115209f
C2426 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 VGND 0.479339f
C2427 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 VGND 0.069002f
C2428 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 VGND 0.2088f
C2429 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 VGND 0.509237f
C2430 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 VGND 0.26045f
C2431 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VGND 0.061029f
C2432 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 VGND 0.019469f
C2433 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 VGND 0.042527f
C2434 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 VGND 0.061029f
C2435 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 VGND 0.019469f
C2436 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 VGND 0.042803f
C2437 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 VGND 0.013718f
C2438 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 VGND 0.061029f
C2439 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VGND 0.019469f
C2440 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 VGND 0.042803f
C2441 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 VGND 0.061029f
C2442 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 VGND 0.019469f
C2443 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 VGND 0.042527f
C2444 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 VGND 0.013568f
C2445 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 VGND 0.358144f
C2446 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 VGND 0.048842f
C2447 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 VGND 0.14784f
C2448 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 VGND 0.375222f
C2449 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 VGND 0.013347f
C2450 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 VGND 0.013347f
C2451 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 VGND 0.031263f
C2452 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 VGND 0.040042f
C2453 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 VGND 0.040042f
C2454 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 VGND 0.081573f
C2455 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 VGND 0.339393f
C2456 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 VGND 0.061913f
C2457 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 VGND 0.061913f
C2458 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 VGND 0.072289f
C2459 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 VGND 0.061913f
C2460 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 VGND 0.061913f
C2461 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 VGND 0.071905f
C2462 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 VGND 0.644548f
C2463 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 VGND 0.046875f
C2464 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 VGND 0.159849f
C2465 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 VGND 0.14784f
C2466 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 VGND 0.245357f
C2467 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 VGND 0.18441f
C2468 a_10958_32492.t5 VGND 0.024913f
C2469 a_10958_32492.t11 VGND 0.096748f
C2470 a_10958_32492.t1 VGND 0.024913f
C2471 a_10958_32492.t12 VGND 0.024913f
C2472 a_10958_32492.n0 VGND 0.060504f
C2473 a_10958_32492.n1 VGND 0.369187f
C2474 a_10958_32492.t10 VGND 0.024913f
C2475 a_10958_32492.t4 VGND 0.024913f
C2476 a_10958_32492.n2 VGND 0.060504f
C2477 a_10958_32492.n3 VGND 0.182084f
C2478 a_10958_32492.t3 VGND 0.024913f
C2479 a_10958_32492.t2 VGND 0.024913f
C2480 a_10958_32492.n4 VGND 0.060504f
C2481 a_10958_32492.n5 VGND 0.221492f
C2482 a_10958_32492.t8 VGND 0.024913f
C2483 a_10958_32492.t0 VGND 0.024913f
C2484 a_10958_32492.n6 VGND 0.052659f
C2485 a_10958_32492.n7 VGND 0.137512f
C2486 a_10958_32492.t6 VGND 0.024913f
C2487 a_10958_32492.t7 VGND 0.024913f
C2488 a_10958_32492.n8 VGND 0.057757f
C2489 a_10958_32492.n9 VGND 0.342225f
C2490 a_10958_32492.n10 VGND 0.059872f
C2491 a_10958_32492.t9 VGND 0.024913f
C2492 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 VGND 0.086195f
C2493 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 VGND 0.027496f
C2494 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 VGND 0.060063f
C2495 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 VGND 0.086195f
C2496 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 VGND 0.027496f
C2497 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 VGND 0.060453f
C2498 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 VGND 0.019374f
C2499 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 VGND 0.086195f
C2500 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 VGND 0.027496f
C2501 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 VGND 0.060453f
C2502 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 VGND 0.086195f
C2503 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 VGND 0.027496f
C2504 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 VGND 0.060063f
C2505 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 VGND 0.019163f
C2506 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 VGND 0.505822f
C2507 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 VGND 0.068982f
C2508 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 VGND 0.2088f
C2509 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 VGND 0.529943f
C2510 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 VGND 0.27612f
C2511 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 VGND 0.018851f
C2512 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 VGND 0.018851f
C2513 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 VGND 0.044154f
C2514 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 VGND 0.056553f
C2515 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 VGND 0.056553f
C2516 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 VGND 0.115209f
C2517 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 VGND 0.479339f
C2518 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 VGND 0.069002f
C2519 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 VGND 0.2088f
C2520 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 VGND 0.509237f
C2521 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 VGND 0.26045f
C2522 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 VGND 0.165681f
C2523 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 VGND 0.051203f
C2524 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 VGND 0.451103f
C2525 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 VGND 0.066664f
C2526 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 VGND 0.021266f
C2527 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 VGND 0.046756f
C2528 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 VGND 0.066664f
C2529 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 VGND 0.021266f
C2530 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 VGND 0.046454f
C2531 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 VGND 0.014982f
C2532 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 VGND 0.066664f
C2533 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 VGND 0.021266f
C2534 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 VGND 0.046756f
C2535 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 VGND 0.066664f
C2536 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 VGND 0.021266f
C2537 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 VGND 0.046454f
C2538 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 VGND 0.014821f
C2539 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 VGND 0.229513f
C2540 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 VGND 0.043739f
C2541 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 VGND 0.043739f
C2542 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 VGND 0.093535f
C2543 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 VGND 0.01458f
C2544 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 VGND 0.01458f
C2545 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 VGND 0.031652f
C2546 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 VGND 0.376142f
C2547 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 VGND 0.165681f
C2548 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 VGND 0.051203f
C2549 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 VGND 0.398173f
C2550 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND 0.027086f
C2551 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VGND 0.034765f
C2552 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VGND 0.034765f
C2553 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 VGND 0.10415f
C2554 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VGND 0.067642f
C2555 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VGND 0.215011f
C2556 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 VGND 0.85898f
C2557 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VGND 0.093153f
C2558 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND 0.086397f
C2559 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VGND 0.093468f
C2560 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 VGND 0.091702f
C2561 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 VGND 0.063806f
C2562 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 VGND 0.942937f
C2563 uo_out[3].t5 VGND 0.007815f
C2564 uo_out[3].t4 VGND 0.026417f
C2565 uo_out[3].n0 VGND 0.021415f
C2566 uo_out[3].t3 VGND 0.015221f
C2567 uo_out[3].t1 VGND 0.015221f
C2568 uo_out[3].n1 VGND 0.032348f
C2569 uo_out[3].n2 VGND 0.141125f
C2570 uo_out[3].t0 VGND 0.005074f
C2571 uo_out[3].t2 VGND 0.005074f
C2572 uo_out[3].n3 VGND 0.011015f
C2573 uo_out[3].n4 VGND 0.037476f
C2574 uo_out[3].n5 VGND 0.713178f
C2575 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 VGND 0.930597f
C2576 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.400887f
C2577 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 VGND 1.11317f
C2578 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.087567f
C2579 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C2580 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.097942f
C2581 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.089004f
C2582 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.08317f
C2583 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C2584 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.041221f
C2585 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.095888f
C2586 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C2587 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.108461f
C2588 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C2589 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C2590 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C2591 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 VGND 0.115417f
C2592 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C2593 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C2594 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.041341f
C2595 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.096169f
C2596 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C2597 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.089265f
C2598 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.083414f
C2599 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C2600 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.202074f
C2601 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C2602 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.03985f
C2603 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C2604 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.200787f
C2605 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C2606 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.054421f
C2607 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C2608 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C2609 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.107523f
C2610 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C2611 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C2612 a_10958_25646.t3 VGND 0.024913f
C2613 a_10958_25646.t4 VGND 0.096748f
C2614 a_10958_25646.t2 VGND 0.024913f
C2615 a_10958_25646.t5 VGND 0.024913f
C2616 a_10958_25646.n0 VGND 0.060504f
C2617 a_10958_25646.n1 VGND 0.369187f
C2618 a_10958_25646.t12 VGND 0.024913f
C2619 a_10958_25646.t1 VGND 0.024913f
C2620 a_10958_25646.n2 VGND 0.060504f
C2621 a_10958_25646.n3 VGND 0.182084f
C2622 a_10958_25646.t0 VGND 0.024913f
C2623 a_10958_25646.t6 VGND 0.024913f
C2624 a_10958_25646.n4 VGND 0.060504f
C2625 a_10958_25646.n5 VGND 0.221492f
C2626 a_10958_25646.t9 VGND 0.024913f
C2627 a_10958_25646.t10 VGND 0.024913f
C2628 a_10958_25646.n6 VGND 0.059872f
C2629 a_10958_25646.t7 VGND 0.024913f
C2630 a_10958_25646.t8 VGND 0.024913f
C2631 a_10958_25646.n7 VGND 0.057757f
C2632 a_10958_25646.n8 VGND 0.342225f
C2633 a_10958_25646.n9 VGND 0.137512f
C2634 a_10958_25646.n10 VGND 0.052659f
C2635 a_10958_25646.t11 VGND 0.024913f
C2636 uo_out[0].t4 VGND 0.012439f
C2637 uo_out[0].t5 VGND 0.042049f
C2638 uo_out[0].n0 VGND 0.034087f
C2639 uo_out[0].t1 VGND 0.024228f
C2640 uo_out[0].t3 VGND 0.024228f
C2641 uo_out[0].n1 VGND 0.051489f
C2642 uo_out[0].n2 VGND 0.224634f
C2643 uo_out[0].t2 VGND 0.008076f
C2644 uo_out[0].t0 VGND 0.008076f
C2645 uo_out[0].n3 VGND 0.017533f
C2646 uo_out[0].n4 VGND 0.059652f
C2647 uo_out[0].n5 VGND 1.71515f
C2648 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 VGND 0.086195f
C2649 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 VGND 0.027496f
C2650 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 VGND 0.060063f
C2651 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 VGND 0.086195f
C2652 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 VGND 0.027496f
C2653 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 VGND 0.060453f
C2654 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 VGND 0.019374f
C2655 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 VGND 0.086195f
C2656 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 VGND 0.027496f
C2657 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 VGND 0.060453f
C2658 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 VGND 0.086195f
C2659 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 VGND 0.027496f
C2660 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 VGND 0.060063f
C2661 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 VGND 0.019163f
C2662 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 VGND 0.505822f
C2663 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 VGND 0.068982f
C2664 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 VGND 0.2088f
C2665 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 VGND 0.529943f
C2666 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 VGND 0.27612f
C2667 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 VGND 0.018851f
C2668 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 VGND 0.018851f
C2669 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 VGND 0.044154f
C2670 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 VGND 0.056553f
C2671 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 VGND 0.056553f
C2672 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 VGND 0.115209f
C2673 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 VGND 0.479339f
C2674 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 VGND 0.069002f
C2675 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 VGND 0.2088f
C2676 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 VGND 0.509237f
C2677 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 VGND 0.26045f
C2678 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 VGND 0.09757f
C2679 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VGND 0.030153f
C2680 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2681 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VGND 0.039259f
C2682 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 VGND 0.012524f
C2683 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2684 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2685 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2686 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2687 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2688 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 VGND 0.039259f
C2689 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2690 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2691 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 VGND 0.039259f
C2692 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2693 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2694 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2695 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2696 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 VGND 0.046129f
C2697 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 VGND 0.046129f
C2698 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2699 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2700 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 VGND 0.046129f
C2701 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2702 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2703 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 VGND 0.025758f
C2704 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 VGND 0.025758f
C2705 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2706 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VGND 0.008586f
C2707 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2708 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2709 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2710 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 VGND 0.09757f
C2711 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 VGND 0.030153f
C2712 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2713 a_10108_30826.t5 VGND 0.059028f
C2714 a_10108_30826.t0 VGND 0.059028f
C2715 a_10108_30826.t3 VGND 0.059028f
C2716 a_10108_30826.n0 VGND 0.136068f
C2717 a_10108_30826.t1 VGND 0.059028f
C2718 a_10108_30826.t2 VGND 0.059028f
C2719 a_10108_30826.n1 VGND 0.258102f
C2720 a_10108_30826.n2 VGND 1.11221f
C2721 a_10108_30826.n3 VGND 0.139449f
C2722 a_10108_30826.t4 VGND 0.059028f
C2723 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 VGND 0.09757f
C2724 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 VGND 0.030153f
C2725 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2726 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VGND 0.039259f
C2727 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 VGND 0.012524f
C2728 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2729 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 VGND 0.039259f
C2730 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2731 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2732 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2733 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2734 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2735 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2736 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 VGND 0.039259f
C2737 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2738 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2739 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2740 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2741 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2742 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 VGND 0.046129f
C2743 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2744 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2745 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 VGND 0.046129f
C2746 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2747 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2748 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 VGND 0.025758f
C2749 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 VGND 0.025758f
C2750 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2751 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2752 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 VGND 0.008586f
C2753 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2754 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2755 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 VGND 0.09757f
C2756 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 VGND 0.030153f
C2757 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2758 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND 0.027086f
C2759 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 VGND 0.034765f
C2760 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 VGND 0.034765f
C2761 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 VGND 0.10415f
C2762 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VGND 0.067642f
C2763 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VGND 0.215011f
C2764 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 VGND 0.85898f
C2765 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND 0.093153f
C2766 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VGND 0.086397f
C2767 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VGND 0.093468f
C2768 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 VGND 0.091702f
C2769 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 VGND 0.063806f
C2770 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 VGND 0.942937f
C2771 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C2772 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C2773 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.087567f
C2774 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C2775 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C2776 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.202442f
C2777 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.089004f
C2778 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C2779 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C2780 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.041221f
C2781 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C2782 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C2783 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C2784 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C2785 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C2786 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.054262f
C2787 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C2788 a_10958_27928.t5 VGND 0.024913f
C2789 a_10958_27928.t4 VGND 0.024913f
C2790 a_10958_27928.t7 VGND 0.024913f
C2791 a_10958_27928.n0 VGND 0.059872f
C2792 a_10958_27928.t3 VGND 0.096748f
C2793 a_10958_27928.t11 VGND 0.024913f
C2794 a_10958_27928.t0 VGND 0.024913f
C2795 a_10958_27928.n1 VGND 0.060504f
C2796 a_10958_27928.n2 VGND 0.369187f
C2797 a_10958_27928.t2 VGND 0.024913f
C2798 a_10958_27928.t9 VGND 0.024913f
C2799 a_10958_27928.n3 VGND 0.060504f
C2800 a_10958_27928.n4 VGND 0.182084f
C2801 a_10958_27928.t12 VGND 0.024913f
C2802 a_10958_27928.t1 VGND 0.024913f
C2803 a_10958_27928.n5 VGND 0.060504f
C2804 a_10958_27928.n6 VGND 0.221492f
C2805 a_10958_27928.t6 VGND 0.024913f
C2806 a_10958_27928.t10 VGND 0.024913f
C2807 a_10958_27928.n7 VGND 0.052659f
C2808 a_10958_27928.n8 VGND 0.137512f
C2809 a_10958_27928.n9 VGND 0.342225f
C2810 a_10958_27928.n10 VGND 0.057757f
C2811 a_10958_27928.t8 VGND 0.024913f
C2812 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 VGND 0.086195f
C2813 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 VGND 0.027496f
C2814 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 VGND 0.060063f
C2815 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 VGND 0.086195f
C2816 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 VGND 0.027496f
C2817 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 VGND 0.060453f
C2818 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 VGND 0.019374f
C2819 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 VGND 0.086195f
C2820 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 VGND 0.027496f
C2821 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 VGND 0.060453f
C2822 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 VGND 0.086195f
C2823 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 VGND 0.027496f
C2824 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 VGND 0.060063f
C2825 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 VGND 0.019163f
C2826 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 VGND 0.505822f
C2827 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 VGND 0.068982f
C2828 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 VGND 0.2088f
C2829 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 VGND 0.529943f
C2830 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 VGND 0.27612f
C2831 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 VGND 0.018851f
C2832 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 VGND 0.018851f
C2833 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 VGND 0.044154f
C2834 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 VGND 0.056553f
C2835 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 VGND 0.056553f
C2836 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 VGND 0.115209f
C2837 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 VGND 0.479339f
C2838 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 VGND 0.069002f
C2839 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 VGND 0.2088f
C2840 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 VGND 0.509237f
C2841 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 VGND 0.26045f
C2842 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 VGND 0.165681f
C2843 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 VGND 0.051203f
C2844 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 VGND 0.451103f
C2845 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 VGND 0.066664f
C2846 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 VGND 0.021266f
C2847 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 VGND 0.046756f
C2848 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 VGND 0.066664f
C2849 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 VGND 0.021266f
C2850 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 VGND 0.046454f
C2851 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 VGND 0.014982f
C2852 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 VGND 0.066664f
C2853 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 VGND 0.021266f
C2854 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 VGND 0.046756f
C2855 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 VGND 0.066664f
C2856 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 VGND 0.021266f
C2857 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 VGND 0.046454f
C2858 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 VGND 0.014821f
C2859 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 VGND 0.229513f
C2860 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 VGND 0.043739f
C2861 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 VGND 0.043739f
C2862 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 VGND 0.093535f
C2863 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 VGND 0.01458f
C2864 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 VGND 0.01458f
C2865 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 VGND 0.031652f
C2866 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 VGND 0.376142f
C2867 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 VGND 0.165681f
C2868 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 VGND 0.051203f
C2869 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 VGND 0.398173f
C2870 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 VGND 0.085944f
C2871 ui_in[5].t5 VGND 0.049226f
C2872 ui_in[5].t7 VGND 0.053255f
C2873 ui_in[5].n0 VGND 0.052248f
C2874 ui_in[5].t3 VGND 0.053075f
C2875 ui_in[5].n1 VGND 0.03636f
C2876 ui_in[5].t4 VGND 0.015432f
C2877 ui_in[5].t6 VGND 0.019808f
C2878 ui_in[5].t2 VGND 0.019808f
C2879 ui_in[5].n2 VGND 0.059369f
C2880 ui_in[5].n3 VGND 0.360373f
C2881 ui_in[5].n4 VGND 2.81694f
C2882 ui_in[5].t0 VGND 0.049902f
C2883 ui_in[5].t1 VGND 0.016108f
C2884 ui_in[5].n5 VGND 0.050487f
C2885 ui_in[5].n6 VGND 0.424074f
C2886 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 VGND 0.019446f
C2887 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 VGND 0.02496f
C2888 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 VGND 0.02496f
C2889 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 VGND 0.074774f
C2890 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 VGND 0.048564f
C2891 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 VGND 0.154367f
C2892 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 VGND 0.616703f
C2893 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 VGND 0.066879f
C2894 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 VGND 0.062029f
C2895 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 VGND 0.067105f
C2896 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 VGND 0.065837f
C2897 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 VGND 0.045809f
C2898 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 VGND 0.676981f
C2899 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 VGND 0.059856f
C2900 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 VGND 0.019094f
C2901 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2902 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 VGND 0.059856f
C2903 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2904 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2905 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2906 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 VGND 0.059856f
C2907 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 VGND 0.019094f
C2908 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2909 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 VGND 0.059856f
C2910 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2911 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2912 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2913 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2914 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 VGND 0.047903f
C2915 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 VGND 0.144997f
C2916 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2917 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 VGND 0.191745f
C2918 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 VGND 0.013091f
C2919 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 VGND 0.013091f
C2920 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 VGND 0.030662f
C2921 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 VGND 0.039272f
C2922 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 VGND 0.039272f
C2923 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 VGND 0.080004f
C2924 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 VGND 0.332866f
C2925 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2926 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 VGND 0.060722f
C2927 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 VGND 0.070899f
C2928 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 VGND 0.060722f
C2929 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 VGND 0.060722f
C2930 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 VGND 0.070523f
C2931 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 VGND 0.632153f
C2932 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 VGND 0.045973f
C2933 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 VGND 0.156775f
C2934 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 VGND 0.144997f
C2935 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 VGND 0.240639f
C2936 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 VGND 0.180864f
C2937 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C2938 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C2939 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.096169f
C2940 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C2941 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C2942 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C2943 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C2944 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C2945 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C2946 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C2947 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.200787f
C2948 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C2949 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.054421f
C2950 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C2951 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C2952 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C2953 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.107523f
C2954 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C2955 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C2956 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VGND 0.09757f
C2957 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VGND 0.030153f
C2958 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2959 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 VGND 0.039259f
C2960 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2961 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2962 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2963 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2964 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2965 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2966 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2967 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2968 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2969 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 VGND 0.039259f
C2970 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 VGND 0.012524f
C2971 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2972 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2973 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2974 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 VGND 0.046129f
C2975 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2976 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2977 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 VGND 0.046129f
C2978 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2979 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2980 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2981 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 VGND 0.025758f
C2982 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 VGND 0.025758f
C2983 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2984 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 VGND 0.008586f
C2985 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 VGND 0.008586f
C2986 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2987 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2988 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 VGND 0.09757f
C2989 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 VGND 0.030153f
C2990 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2991 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 VGND 0.165681f
C2992 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 VGND 0.051203f
C2993 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 VGND 0.451103f
C2994 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 VGND 0.066664f
C2995 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 VGND 0.021266f
C2996 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 VGND 0.046756f
C2997 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 VGND 0.066664f
C2998 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 VGND 0.021266f
C2999 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 VGND 0.046454f
C3000 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 VGND 0.014982f
C3001 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 VGND 0.066664f
C3002 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 VGND 0.021266f
C3003 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 VGND 0.046756f
C3004 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 VGND 0.066664f
C3005 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 VGND 0.021266f
C3006 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 VGND 0.046454f
C3007 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 VGND 0.014821f
C3008 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 VGND 0.229513f
C3009 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 VGND 0.043739f
C3010 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 VGND 0.043739f
C3011 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 VGND 0.093535f
C3012 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 VGND 0.01458f
C3013 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 VGND 0.01458f
C3014 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 VGND 0.031652f
C3015 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 VGND 0.376142f
C3016 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 VGND 0.165681f
C3017 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 VGND 0.051203f
C3018 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 VGND 0.398173f
C3019 a_10958_34774.t4 VGND 0.024913f
C3020 a_10958_34774.t5 VGND 0.024913f
C3021 a_10958_34774.t7 VGND 0.024913f
C3022 a_10958_34774.n0 VGND 0.059872f
C3023 a_10958_34774.t12 VGND 0.096748f
C3024 a_10958_34774.t11 VGND 0.024913f
C3025 a_10958_34774.t2 VGND 0.024913f
C3026 a_10958_34774.n1 VGND 0.060504f
C3027 a_10958_34774.n2 VGND 0.369187f
C3028 a_10958_34774.t1 VGND 0.024913f
C3029 a_10958_34774.t10 VGND 0.024913f
C3030 a_10958_34774.n3 VGND 0.060504f
C3031 a_10958_34774.n4 VGND 0.182084f
C3032 a_10958_34774.t3 VGND 0.024913f
C3033 a_10958_34774.t0 VGND 0.024913f
C3034 a_10958_34774.n5 VGND 0.060504f
C3035 a_10958_34774.n6 VGND 0.221492f
C3036 a_10958_34774.t6 VGND 0.024913f
C3037 a_10958_34774.t9 VGND 0.024913f
C3038 a_10958_34774.n7 VGND 0.052659f
C3039 a_10958_34774.n8 VGND 0.137512f
C3040 a_10958_34774.n9 VGND 0.342225f
C3041 a_10958_34774.n10 VGND 0.057757f
C3042 a_10958_34774.t8 VGND 0.024913f
C3043 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 VGND 0.060722f
C3044 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 VGND 0.060722f
C3045 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 VGND 0.070899f
C3046 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 VGND 0.060722f
C3047 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 VGND 0.060722f
C3048 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 VGND 0.070523f
C3049 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 VGND 0.632153f
C3050 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 VGND 0.059856f
C3051 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 VGND 0.019094f
C3052 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 VGND 0.041709f
C3053 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 VGND 0.059856f
C3054 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 VGND 0.019094f
C3055 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 VGND 0.04198f
C3056 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 VGND 0.013454f
C3057 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VGND 0.059856f
C3058 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VGND 0.019094f
C3059 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 VGND 0.04198f
C3060 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 VGND 0.059856f
C3061 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 VGND 0.019094f
C3062 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 VGND 0.041709f
C3063 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 VGND 0.013307f
C3064 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 VGND 0.351257f
C3065 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 VGND 0.047903f
C3066 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VGND 0.144997f
C3067 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 VGND 0.368007f
C3068 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VGND 0.013091f
C3069 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 VGND 0.013091f
C3070 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 VGND 0.030662f
C3071 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 VGND 0.039272f
C3072 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 VGND 0.039272f
C3073 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 VGND 0.080004f
C3074 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 VGND 0.332866f
C3075 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 VGND 0.180864f
C3076 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 VGND 0.144997f
C3077 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 VGND 0.240639f
C3078 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 VGND 0.045973f
C3079 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 VGND 0.156775f
C3080 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 VGND 0.086195f
C3081 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 VGND 0.027496f
C3082 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 VGND 0.060063f
C3083 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 VGND 0.086195f
C3084 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 VGND 0.027496f
C3085 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 VGND 0.060453f
C3086 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 VGND 0.019374f
C3087 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 VGND 0.086195f
C3088 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 VGND 0.027496f
C3089 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 VGND 0.060453f
C3090 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 VGND 0.086195f
C3091 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 VGND 0.027496f
C3092 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 VGND 0.060063f
C3093 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 VGND 0.019163f
C3094 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 VGND 0.505822f
C3095 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 VGND 0.068982f
C3096 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 VGND 0.2088f
C3097 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 VGND 0.529943f
C3098 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 VGND 0.302329f
C3099 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 VGND 0.018851f
C3100 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 VGND 0.018851f
C3101 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 VGND 0.044154f
C3102 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 VGND 0.056553f
C3103 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 VGND 0.056553f
C3104 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 VGND 0.115209f
C3105 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 VGND 0.479339f
C3106 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 VGND 0.069002f
C3107 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 VGND 0.2088f
C3108 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 VGND 0.509237f
C3109 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 VGND 0.26045f
C3110 tdc_0.diff_gen_0.delay_unit_2_4.out_1 VGND 0.212791f
C3111 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 VGND 0.165681f
C3112 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 VGND 0.051203f
C3113 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 VGND 0.451103f
C3114 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 VGND 0.066664f
C3115 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 VGND 0.021266f
C3116 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 VGND 0.046756f
C3117 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 VGND 0.066664f
C3118 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 VGND 0.021266f
C3119 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 VGND 0.046454f
C3120 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 VGND 0.014982f
C3121 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 VGND 0.066664f
C3122 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 VGND 0.021266f
C3123 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 VGND 0.046756f
C3124 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 VGND 0.066664f
C3125 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 VGND 0.021266f
C3126 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 VGND 0.046454f
C3127 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 VGND 0.014821f
C3128 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 VGND 0.229513f
C3129 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 VGND 0.043739f
C3130 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 VGND 0.043739f
C3131 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 VGND 0.093535f
C3132 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 VGND 0.01458f
C3133 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 VGND 0.01458f
C3134 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 VGND 0.031652f
C3135 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 VGND 0.376142f
C3136 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 VGND 0.165681f
C3137 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 VGND 0.051203f
C3138 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 VGND 0.398173f
C3139 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 VGND 0.086195f
C3140 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 VGND 0.027496f
C3141 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 VGND 0.060063f
C3142 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 VGND 0.086195f
C3143 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 VGND 0.027496f
C3144 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 VGND 0.060453f
C3145 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 VGND 0.019374f
C3146 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 VGND 0.086195f
C3147 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 VGND 0.027496f
C3148 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 VGND 0.060453f
C3149 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 VGND 0.086195f
C3150 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 VGND 0.027496f
C3151 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 VGND 0.060063f
C3152 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 VGND 0.019163f
C3153 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 VGND 0.505822f
C3154 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 VGND 0.068982f
C3155 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 VGND 0.2088f
C3156 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 VGND 0.529943f
C3157 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 VGND 0.27612f
C3158 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 VGND 0.018851f
C3159 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 VGND 0.018851f
C3160 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 VGND 0.044154f
C3161 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 VGND 0.056553f
C3162 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 VGND 0.056553f
C3163 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 VGND 0.115209f
C3164 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 VGND 0.479339f
C3165 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 VGND 0.069002f
C3166 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 VGND 0.2088f
C3167 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 VGND 0.509237f
C3168 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 VGND 0.26045f
C3169 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 VGND 0.165681f
C3170 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 VGND 0.051203f
C3171 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 VGND 0.451103f
C3172 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 VGND 0.066664f
C3173 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 VGND 0.021266f
C3174 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 VGND 0.046756f
C3175 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 VGND 0.066664f
C3176 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 VGND 0.021266f
C3177 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 VGND 0.046454f
C3178 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 VGND 0.014982f
C3179 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 VGND 0.066664f
C3180 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 VGND 0.021266f
C3181 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 VGND 0.046756f
C3182 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 VGND 0.066664f
C3183 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 VGND 0.021266f
C3184 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 VGND 0.046454f
C3185 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 VGND 0.014821f
C3186 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 VGND 0.229513f
C3187 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 VGND 0.043739f
C3188 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 VGND 0.043739f
C3189 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 VGND 0.093535f
C3190 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 VGND 0.01458f
C3191 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 VGND 0.01458f
C3192 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 VGND 0.031652f
C3193 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 VGND 0.376142f
C3194 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 VGND 0.165681f
C3195 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 VGND 0.051203f
C3196 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 VGND 0.398173f
C3197 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 VGND 0.085944f
C3198 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 VGND 0.019446f
C3199 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 VGND 0.02496f
C3200 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 VGND 0.02496f
C3201 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 VGND 0.074774f
C3202 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 VGND 0.048564f
C3203 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 VGND 0.154367f
C3204 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 VGND 0.616703f
C3205 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 VGND 0.066879f
C3206 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 VGND 0.062029f
C3207 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 VGND 0.067105f
C3208 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 VGND 0.065837f
C3209 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 VGND 0.045809f
C3210 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 VGND 0.676981f
C3211 a_10108_26262.t1 VGND 0.059028f
C3212 a_10108_26262.t3 VGND 0.059028f
C3213 a_10108_26262.t5 VGND 0.059028f
C3214 a_10108_26262.n0 VGND 0.136068f
C3215 a_10108_26262.t4 VGND 0.059028f
C3216 a_10108_26262.t0 VGND 0.059028f
C3217 a_10108_26262.n1 VGND 0.258102f
C3218 a_10108_26262.n2 VGND 1.11221f
C3219 a_10108_26262.n3 VGND 0.139449f
C3220 a_10108_26262.t2 VGND 0.059028f
C3221 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3222 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.041341f
C3223 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.096169f
C3224 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3225 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.089265f
C3226 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.083414f
C3227 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3228 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C3229 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.03985f
C3230 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3231 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C3232 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.202074f
C3233 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C3234 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3235 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3236 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3237 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.107523f
C3238 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3239 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3240 a_10958_37056.t6 VGND 0.024913f
C3241 a_10958_37056.t7 VGND 0.024913f
C3242 a_10958_37056.t4 VGND 0.024913f
C3243 a_10958_37056.n0 VGND 0.059872f
C3244 a_10958_37056.t11 VGND 0.096748f
C3245 a_10958_37056.t0 VGND 0.024913f
C3246 a_10958_37056.t10 VGND 0.024913f
C3247 a_10958_37056.n1 VGND 0.060504f
C3248 a_10958_37056.n2 VGND 0.369187f
C3249 a_10958_37056.t12 VGND 0.024913f
C3250 a_10958_37056.t1 VGND 0.024913f
C3251 a_10958_37056.n3 VGND 0.060504f
C3252 a_10958_37056.n4 VGND 0.182084f
C3253 a_10958_37056.t9 VGND 0.024913f
C3254 a_10958_37056.t2 VGND 0.024913f
C3255 a_10958_37056.n5 VGND 0.060504f
C3256 a_10958_37056.n6 VGND 0.221492f
C3257 a_10958_37056.t5 VGND 0.024913f
C3258 a_10958_37056.t3 VGND 0.024913f
C3259 a_10958_37056.n7 VGND 0.052659f
C3260 a_10958_37056.n8 VGND 0.137512f
C3261 a_10958_37056.n9 VGND 0.342225f
C3262 a_10958_37056.n10 VGND 0.057757f
C3263 a_10958_37056.t8 VGND 0.024913f
C3264 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 VGND 0.027086f
C3265 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 VGND 0.034765f
C3266 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 VGND 0.034765f
C3267 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 VGND 0.10415f
C3268 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 VGND 0.067642f
C3269 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 VGND 0.215011f
C3270 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 VGND 0.85898f
C3271 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 VGND 0.093153f
C3272 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 VGND 0.086397f
C3273 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 VGND 0.093468f
C3274 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 VGND 0.091702f
C3275 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 VGND 0.063806f
C3276 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 VGND 0.942937f
C3277 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 VGND 0.375772f
C3278 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d VGND 0.696742f
C3279 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 VGND 0.059856f
C3280 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 VGND 0.019094f
C3281 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 VGND 0.041709f
C3282 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 VGND 0.059856f
C3283 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 VGND 0.019094f
C3284 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 VGND 0.04198f
C3285 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 VGND 0.013454f
C3286 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VGND 0.059856f
C3287 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VGND 0.019094f
C3288 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 VGND 0.04198f
C3289 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 VGND 0.059856f
C3290 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 VGND 0.019094f
C3291 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 VGND 0.041709f
C3292 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 VGND 0.013307f
C3293 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 VGND 0.351257f
C3294 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 VGND 0.047903f
C3295 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 VGND 0.144997f
C3296 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 VGND 0.368007f
C3297 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 VGND 0.013091f
C3298 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 VGND 0.013091f
C3299 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 VGND 0.030662f
C3300 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 VGND 0.039272f
C3301 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 VGND 0.039272f
C3302 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 VGND 0.080004f
C3303 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 VGND 0.332866f
C3304 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 VGND 0.060722f
C3305 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 VGND 0.060722f
C3306 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 VGND 0.070899f
C3307 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 VGND 0.060722f
C3308 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 VGND 0.060722f
C3309 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 VGND 0.070523f
C3310 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 VGND 0.632153f
C3311 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 VGND 0.045973f
C3312 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 VGND 0.156775f
C3313 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 VGND 0.144997f
C3314 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 VGND 0.240639f
C3315 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 VGND 0.180864f
C3316 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 VGND 0.271416f
C3317 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 VGND 0.019446f
C3318 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 VGND 0.02496f
C3319 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 VGND 0.02496f
C3320 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 VGND 0.074774f
C3321 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 VGND 0.048564f
C3322 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 VGND 0.154367f
C3323 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 VGND 0.616703f
C3324 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 VGND 0.066879f
C3325 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 VGND 0.062029f
C3326 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 VGND 0.067105f
C3327 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 VGND 0.065837f
C3328 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 VGND 0.045809f
C3329 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 VGND 0.676981f
C3330 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3331 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3332 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3333 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3334 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.089265f
C3335 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3336 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3337 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C3338 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C3339 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.03985f
C3340 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3341 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C3342 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3343 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3344 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3345 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3346 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C3347 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3348 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3349 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3350 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3351 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.087567f
C3352 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.039734f
C3353 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3354 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.089004f
C3355 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.08317f
C3356 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C3357 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.041221f
C3358 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C3359 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C3360 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.108461f
C3361 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C3362 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3363 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.054262f
C3364 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C3365 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3366 a_10108_35390.t1 VGND 0.059028f
C3367 a_10108_35390.t3 VGND 0.059028f
C3368 a_10108_35390.t0 VGND 0.059028f
C3369 a_10108_35390.n0 VGND 0.136068f
C3370 a_10108_35390.t4 VGND 0.059028f
C3371 a_10108_35390.t5 VGND 0.059028f
C3372 a_10108_35390.n1 VGND 0.258102f
C3373 a_10108_35390.n2 VGND 1.11221f
C3374 a_10108_35390.n3 VGND 0.139449f
C3375 a_10108_35390.t2 VGND 0.059028f
C3376 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3377 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3378 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.087567f
C3379 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.039734f
C3380 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3381 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C3382 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.089004f
C3383 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.08317f
C3384 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C3385 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.041221f
C3386 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.095888f
C3387 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C3388 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.108461f
C3389 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C3390 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.054262f
C3391 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3392 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C3393 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3394 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3395 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3396 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3397 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.089265f
C3398 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3399 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3400 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.087824f
C3401 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3402 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3403 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C3404 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C3405 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3406 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3407 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3408 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3409 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.107523f
C3410 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3411 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3412 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3413 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3414 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.087567f
C3415 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.039734f
C3416 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3417 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.089004f
C3418 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.08317f
C3419 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C3420 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.041221f
C3421 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C3422 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C3423 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.108461f
C3424 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.202442f
C3425 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C3426 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.054262f
C3427 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C3428 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3429 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND 0.019446f
C3430 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VGND 0.02496f
C3431 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VGND 0.02496f
C3432 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 VGND 0.074774f
C3433 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VGND 0.048564f
C3434 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VGND 0.154367f
C3435 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 VGND 0.616703f
C3436 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VGND 0.066879f
C3437 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND 0.062029f
C3438 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VGND 0.067105f
C3439 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 VGND 0.065837f
C3440 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 VGND 0.045809f
C3441 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 VGND 0.676981f
C3442 a_10958_23364.t6 VGND 0.024913f
C3443 a_10958_23364.t1 VGND 0.096748f
C3444 a_10958_23364.t9 VGND 0.024913f
C3445 a_10958_23364.t2 VGND 0.024913f
C3446 a_10958_23364.n0 VGND 0.060504f
C3447 a_10958_23364.n1 VGND 0.369187f
C3448 a_10958_23364.t0 VGND 0.024913f
C3449 a_10958_23364.t10 VGND 0.024913f
C3450 a_10958_23364.n2 VGND 0.060504f
C3451 a_10958_23364.n3 VGND 0.182084f
C3452 a_10958_23364.t12 VGND 0.024913f
C3453 a_10958_23364.t8 VGND 0.024913f
C3454 a_10958_23364.n4 VGND 0.060504f
C3455 a_10958_23364.n5 VGND 0.221492f
C3456 a_10958_23364.t3 VGND 0.024913f
C3457 a_10958_23364.t11 VGND 0.024913f
C3458 a_10958_23364.n6 VGND 0.052659f
C3459 a_10958_23364.n7 VGND 0.137512f
C3460 a_10958_23364.t4 VGND 0.024913f
C3461 a_10958_23364.t5 VGND 0.024913f
C3462 a_10958_23364.n8 VGND 0.057757f
C3463 a_10958_23364.n9 VGND 0.342225f
C3464 a_10958_23364.n10 VGND 0.059872f
C3465 a_10958_23364.t7 VGND 0.024913f
C3466 a_10108_28544.t0 VGND 0.059028f
C3467 a_10108_28544.t5 VGND 0.059028f
C3468 a_10108_28544.t2 VGND 0.059028f
C3469 a_10108_28544.n0 VGND 0.136068f
C3470 a_10108_28544.t3 VGND 0.059028f
C3471 a_10108_28544.t4 VGND 0.059028f
C3472 a_10108_28544.n1 VGND 0.258102f
C3473 a_10108_28544.n2 VGND 1.11221f
C3474 a_10108_28544.n3 VGND 0.139449f
C3475 a_10108_28544.t1 VGND 0.059028f
C3476 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3477 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3478 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.087567f
C3479 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C3480 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3481 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C3482 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3483 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C3484 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C3485 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.089004f
C3486 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C3487 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C3488 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C3489 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C3490 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C3491 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.108461f
C3492 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3493 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3494 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3495 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.096169f
C3496 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3497 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C3498 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3499 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3500 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C3501 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3502 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3503 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C3504 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C3505 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3506 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3507 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3508 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3509 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C3510 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3511 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3512 a_10958_39338.t4 VGND 0.024913f
C3513 a_10958_39338.t0 VGND 0.096748f
C3514 a_10958_39338.t8 VGND 0.024913f
C3515 a_10958_39338.t2 VGND 0.024913f
C3516 a_10958_39338.n0 VGND 0.060504f
C3517 a_10958_39338.n1 VGND 0.369187f
C3518 a_10958_39338.t1 VGND 0.024913f
C3519 a_10958_39338.t11 VGND 0.024913f
C3520 a_10958_39338.n2 VGND 0.060504f
C3521 a_10958_39338.n3 VGND 0.182084f
C3522 a_10958_39338.t9 VGND 0.024913f
C3523 a_10958_39338.t12 VGND 0.024913f
C3524 a_10958_39338.n4 VGND 0.060504f
C3525 a_10958_39338.n5 VGND 0.221492f
C3526 a_10958_39338.t3 VGND 0.024913f
C3527 a_10958_39338.t10 VGND 0.024913f
C3528 a_10958_39338.n6 VGND 0.052659f
C3529 a_10958_39338.n7 VGND 0.137512f
C3530 a_10958_39338.t5 VGND 0.024913f
C3531 a_10958_39338.t6 VGND 0.024913f
C3532 a_10958_39338.n8 VGND 0.057757f
C3533 a_10958_39338.n9 VGND 0.342225f
C3534 a_10958_39338.n10 VGND 0.059872f
C3535 a_10958_39338.t7 VGND 0.024913f
C3536 a_10108_39954.t1 VGND 0.059028f
C3537 a_10108_39954.t3 VGND 0.059028f
C3538 a_10108_39954.t2 VGND 0.059028f
C3539 a_10108_39954.n0 VGND 0.136068f
C3540 a_10108_39954.t4 VGND 0.059028f
C3541 a_10108_39954.t5 VGND 0.059028f
C3542 a_10108_39954.n1 VGND 0.258102f
C3543 a_10108_39954.n2 VGND 1.11221f
C3544 a_10108_39954.n3 VGND 0.139449f
C3545 a_10108_39954.t0 VGND 0.059028f
C3546 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd VGND 0.503525f
C3547 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 VGND 0.130197f
C3548 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 VGND 0.189073f
C3549 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 VGND 0.025758f
C3550 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 VGND 0.025758f
C3551 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 VGND 0.055083f
C3552 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 VGND 0.008586f
C3553 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 VGND 0.008586f
C3554 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 VGND 0.01864f
C3555 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 VGND 0.221512f
C3556 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 VGND 0.09757f
C3557 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 VGND 0.030153f
C3558 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 VGND 0.234486f
C3559 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 VGND 0.046129f
C3560 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 VGND 0.046129f
C3561 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 VGND 0.054044f
C3562 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 VGND 0.046129f
C3563 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 VGND 0.046129f
C3564 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 VGND 0.0538f
C3565 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 VGND 0.495704f
C3566 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VGND 0.09757f
C3567 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VGND 0.030153f
C3568 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 VGND 0.265657f
C3569 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 VGND 0.039259f
C3570 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 VGND 0.012524f
C3571 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 VGND 0.027534f
C3572 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 VGND 0.039259f
C3573 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 VGND 0.012524f
C3574 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 VGND 0.027357f
C3575 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 VGND 0.008823f
C3576 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 VGND 0.039259f
C3577 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 VGND 0.012524f
C3578 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 VGND 0.027534f
C3579 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 VGND 0.039259f
C3580 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 VGND 0.012524f
C3581 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 VGND 0.027357f
C3582 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 VGND 0.008728f
C3583 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 VGND 0.135162f
C3584 tdc_0.vernier_delay_line_0.stop_strong.t78 VGND 0.078403f
C3585 tdc_0.vernier_delay_line_0.stop_strong.t43 VGND 0.073263f
C3586 tdc_0.vernier_delay_line_0.stop_strong.n0 VGND 0.070349f
C3587 tdc_0.vernier_delay_line_0.stop_strong.t55 VGND 0.073263f
C3588 tdc_0.vernier_delay_line_0.stop_strong.n1 VGND 0.040134f
C3589 tdc_0.vernier_delay_line_0.stop_strong.t72 VGND 0.073263f
C3590 tdc_0.vernier_delay_line_0.stop_strong.n2 VGND 0.040134f
C3591 tdc_0.vernier_delay_line_0.stop_strong.t37 VGND 0.073263f
C3592 tdc_0.vernier_delay_line_0.stop_strong.n3 VGND 0.064514f
C3593 tdc_0.vernier_delay_line_0.stop_strong.t56 VGND 0.093756f
C3594 tdc_0.vernier_delay_line_0.stop_strong.t87 VGND 0.093545f
C3595 tdc_0.vernier_delay_line_0.stop_strong.n4 VGND 0.403473f
C3596 tdc_0.vernier_delay_line_0.stop_strong.n5 VGND 0.933667f
C3597 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk VGND 1.3151f
C3598 tdc_0.vernier_delay_line_0.stop_strong.t67 VGND 0.078403f
C3599 tdc_0.vernier_delay_line_0.stop_strong.t33 VGND 0.073263f
C3600 tdc_0.vernier_delay_line_0.stop_strong.n6 VGND 0.070349f
C3601 tdc_0.vernier_delay_line_0.stop_strong.t60 VGND 0.073263f
C3602 tdc_0.vernier_delay_line_0.stop_strong.n7 VGND 0.040134f
C3603 tdc_0.vernier_delay_line_0.stop_strong.t82 VGND 0.073263f
C3604 tdc_0.vernier_delay_line_0.stop_strong.n8 VGND 0.040134f
C3605 tdc_0.vernier_delay_line_0.stop_strong.t46 VGND 0.073263f
C3606 tdc_0.vernier_delay_line_0.stop_strong.n9 VGND 0.064514f
C3607 tdc_0.vernier_delay_line_0.stop_strong.t80 VGND 0.093756f
C3608 tdc_0.vernier_delay_line_0.stop_strong.t39 VGND 0.093545f
C3609 tdc_0.vernier_delay_line_0.stop_strong.n10 VGND 0.403473f
C3610 tdc_0.vernier_delay_line_0.stop_strong.n11 VGND 0.777822f
C3611 tdc_0.vernier_delay_line_0.stop_strong.n12 VGND 0.697925f
C3612 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3613 tdc_0.vernier_delay_line_0.stop_strong.t52 VGND 0.078403f
C3614 tdc_0.vernier_delay_line_0.stop_strong.t68 VGND 0.073263f
C3615 tdc_0.vernier_delay_line_0.stop_strong.n13 VGND 0.070349f
C3616 tdc_0.vernier_delay_line_0.stop_strong.t35 VGND 0.073263f
C3617 tdc_0.vernier_delay_line_0.stop_strong.n14 VGND 0.040134f
C3618 tdc_0.vernier_delay_line_0.stop_strong.t51 VGND 0.073263f
C3619 tdc_0.vernier_delay_line_0.stop_strong.n15 VGND 0.040134f
C3620 tdc_0.vernier_delay_line_0.stop_strong.t64 VGND 0.073263f
C3621 tdc_0.vernier_delay_line_0.stop_strong.n16 VGND 0.064514f
C3622 tdc_0.vernier_delay_line_0.stop_strong.t61 VGND 0.093756f
C3623 tdc_0.vernier_delay_line_0.stop_strong.t59 VGND 0.093545f
C3624 tdc_0.vernier_delay_line_0.stop_strong.n17 VGND 0.403473f
C3625 tdc_0.vernier_delay_line_0.stop_strong.n18 VGND 0.777822f
C3626 tdc_0.vernier_delay_line_0.stop_strong.n19 VGND 0.697925f
C3627 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3628 tdc_0.vernier_delay_line_0.stop_strong.t40 VGND 0.078403f
C3629 tdc_0.vernier_delay_line_0.stop_strong.t53 VGND 0.073263f
C3630 tdc_0.vernier_delay_line_0.stop_strong.n20 VGND 0.070349f
C3631 tdc_0.vernier_delay_line_0.stop_strong.t69 VGND 0.073263f
C3632 tdc_0.vernier_delay_line_0.stop_strong.n21 VGND 0.040134f
C3633 tdc_0.vernier_delay_line_0.stop_strong.t71 VGND 0.073263f
C3634 tdc_0.vernier_delay_line_0.stop_strong.n22 VGND 0.040134f
C3635 tdc_0.vernier_delay_line_0.stop_strong.t36 VGND 0.073263f
C3636 tdc_0.vernier_delay_line_0.stop_strong.n23 VGND 0.064514f
C3637 tdc_0.vernier_delay_line_0.stop_strong.t49 VGND 0.093756f
C3638 tdc_0.vernier_delay_line_0.stop_strong.t45 VGND 0.093545f
C3639 tdc_0.vernier_delay_line_0.stop_strong.n24 VGND 0.403473f
C3640 tdc_0.vernier_delay_line_0.stop_strong.n25 VGND 0.777822f
C3641 tdc_0.vernier_delay_line_0.stop_strong.n26 VGND 0.697925f
C3642 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3643 tdc_0.vernier_delay_line_0.stop_strong.t70 VGND 0.078403f
C3644 tdc_0.vernier_delay_line_0.stop_strong.t42 VGND 0.073263f
C3645 tdc_0.vernier_delay_line_0.stop_strong.n27 VGND 0.070349f
C3646 tdc_0.vernier_delay_line_0.stop_strong.t44 VGND 0.073263f
C3647 tdc_0.vernier_delay_line_0.stop_strong.n28 VGND 0.040134f
C3648 tdc_0.vernier_delay_line_0.stop_strong.t57 VGND 0.073263f
C3649 tdc_0.vernier_delay_line_0.stop_strong.n29 VGND 0.040134f
C3650 tdc_0.vernier_delay_line_0.stop_strong.t73 VGND 0.073263f
C3651 tdc_0.vernier_delay_line_0.stop_strong.n30 VGND 0.064514f
C3652 tdc_0.vernier_delay_line_0.stop_strong.t66 VGND 0.093756f
C3653 tdc_0.vernier_delay_line_0.stop_strong.t77 VGND 0.093545f
C3654 tdc_0.vernier_delay_line_0.stop_strong.n31 VGND 0.403473f
C3655 tdc_0.vernier_delay_line_0.stop_strong.n32 VGND 0.777822f
C3656 tdc_0.vernier_delay_line_0.stop_strong.n33 VGND 0.697925f
C3657 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3658 tdc_0.vernier_delay_line_0.stop_strong.t81 VGND 0.078403f
C3659 tdc_0.vernier_delay_line_0.stop_strong.t83 VGND 0.073263f
C3660 tdc_0.vernier_delay_line_0.stop_strong.n34 VGND 0.070349f
C3661 tdc_0.vernier_delay_line_0.stop_strong.t47 VGND 0.073263f
C3662 tdc_0.vernier_delay_line_0.stop_strong.n35 VGND 0.040134f
C3663 tdc_0.vernier_delay_line_0.stop_strong.t62 VGND 0.073263f
C3664 tdc_0.vernier_delay_line_0.stop_strong.n36 VGND 0.040134f
C3665 tdc_0.vernier_delay_line_0.stop_strong.t84 VGND 0.073263f
C3666 tdc_0.vernier_delay_line_0.stop_strong.n37 VGND 0.064514f
C3667 tdc_0.vernier_delay_line_0.stop_strong.t76 VGND 0.093756f
C3668 tdc_0.vernier_delay_line_0.stop_strong.t74 VGND 0.093545f
C3669 tdc_0.vernier_delay_line_0.stop_strong.n38 VGND 0.403473f
C3670 tdc_0.vernier_delay_line_0.stop_strong.n39 VGND 0.777822f
C3671 tdc_0.vernier_delay_line_0.stop_strong.n40 VGND 0.697925f
C3672 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3673 tdc_0.vernier_delay_line_0.stop_strong.t38 VGND 0.078403f
C3674 tdc_0.vernier_delay_line_0.stop_strong.t65 VGND 0.073263f
C3675 tdc_0.vernier_delay_line_0.stop_strong.n41 VGND 0.070349f
C3676 tdc_0.vernier_delay_line_0.stop_strong.t85 VGND 0.073263f
C3677 tdc_0.vernier_delay_line_0.stop_strong.n42 VGND 0.040134f
C3678 tdc_0.vernier_delay_line_0.stop_strong.t50 VGND 0.073263f
C3679 tdc_0.vernier_delay_line_0.stop_strong.n43 VGND 0.040134f
C3680 tdc_0.vernier_delay_line_0.stop_strong.t63 VGND 0.073263f
C3681 tdc_0.vernier_delay_line_0.stop_strong.n44 VGND 0.064514f
C3682 tdc_0.vernier_delay_line_0.stop_strong.t48 VGND 0.093756f
C3683 tdc_0.vernier_delay_line_0.stop_strong.t58 VGND 0.093545f
C3684 tdc_0.vernier_delay_line_0.stop_strong.n45 VGND 0.403473f
C3685 tdc_0.vernier_delay_line_0.stop_strong.n46 VGND 0.777822f
C3686 tdc_0.vernier_delay_line_0.stop_strong.n47 VGND 0.697925f
C3687 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3688 tdc_0.vernier_delay_line_0.stop_strong.t75 VGND 0.078403f
C3689 tdc_0.vernier_delay_line_0.stop_strong.t41 VGND 0.073263f
C3690 tdc_0.vernier_delay_line_0.stop_strong.n48 VGND 0.070349f
C3691 tdc_0.vernier_delay_line_0.stop_strong.t54 VGND 0.073263f
C3692 tdc_0.vernier_delay_line_0.stop_strong.n49 VGND 0.040134f
C3693 tdc_0.vernier_delay_line_0.stop_strong.t32 VGND 0.073263f
C3694 tdc_0.vernier_delay_line_0.stop_strong.n50 VGND 0.040134f
C3695 tdc_0.vernier_delay_line_0.stop_strong.t34 VGND 0.073263f
C3696 tdc_0.vernier_delay_line_0.stop_strong.n51 VGND 0.064514f
C3697 tdc_0.vernier_delay_line_0.stop_strong.t86 VGND 0.093756f
C3698 tdc_0.vernier_delay_line_0.stop_strong.t79 VGND 0.093545f
C3699 tdc_0.vernier_delay_line_0.stop_strong.n52 VGND 0.403473f
C3700 tdc_0.vernier_delay_line_0.stop_strong.n53 VGND 0.777822f
C3701 tdc_0.vernier_delay_line_0.stop_strong.n54 VGND 0.697925f
C3702 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk VGND 0.971005f
C3703 tdc_0.vernier_delay_line_0.stop_strong.t27 VGND 0.181057f
C3704 tdc_0.vernier_delay_line_0.stop_strong.t13 VGND 0.055955f
C3705 tdc_0.vernier_delay_line_0.stop_strong.n55 VGND 0.420822f
C3706 tdc_0.vernier_delay_line_0.stop_strong.t20 VGND 0.181057f
C3707 tdc_0.vernier_delay_line_0.stop_strong.t6 VGND 0.055955f
C3708 tdc_0.vernier_delay_line_0.stop_strong.n56 VGND 0.413796f
C3709 tdc_0.vernier_delay_line_0.stop_strong.n57 VGND 0.17535f
C3710 tdc_0.vernier_delay_line_0.stop_strong.t30 VGND 0.181057f
C3711 tdc_0.vernier_delay_line_0.stop_strong.t0 VGND 0.055955f
C3712 tdc_0.vernier_delay_line_0.stop_strong.n58 VGND 0.413796f
C3713 tdc_0.vernier_delay_line_0.stop_strong.n59 VGND 0.11234f
C3714 tdc_0.vernier_delay_line_0.stop_strong.t23 VGND 0.181057f
C3715 tdc_0.vernier_delay_line_0.stop_strong.t9 VGND 0.055955f
C3716 tdc_0.vernier_delay_line_0.stop_strong.n60 VGND 0.413796f
C3717 tdc_0.vernier_delay_line_0.stop_strong.n61 VGND 0.11234f
C3718 tdc_0.vernier_delay_line_0.stop_strong.t17 VGND 0.181057f
C3719 tdc_0.vernier_delay_line_0.stop_strong.t3 VGND 0.055955f
C3720 tdc_0.vernier_delay_line_0.stop_strong.n62 VGND 0.413796f
C3721 tdc_0.vernier_delay_line_0.stop_strong.n63 VGND 0.11234f
C3722 tdc_0.vernier_delay_line_0.stop_strong.t26 VGND 0.181057f
C3723 tdc_0.vernier_delay_line_0.stop_strong.t12 VGND 0.055955f
C3724 tdc_0.vernier_delay_line_0.stop_strong.n64 VGND 0.413796f
C3725 tdc_0.vernier_delay_line_0.stop_strong.n65 VGND 0.11234f
C3726 tdc_0.vernier_delay_line_0.stop_strong.t16 VGND 0.181057f
C3727 tdc_0.vernier_delay_line_0.stop_strong.t2 VGND 0.055955f
C3728 tdc_0.vernier_delay_line_0.stop_strong.n66 VGND 0.413796f
C3729 tdc_0.vernier_delay_line_0.stop_strong.n67 VGND 0.11234f
C3730 tdc_0.vernier_delay_line_0.stop_strong.t25 VGND 0.181057f
C3731 tdc_0.vernier_delay_line_0.stop_strong.t11 VGND 0.055955f
C3732 tdc_0.vernier_delay_line_0.stop_strong.n68 VGND 0.413796f
C3733 tdc_0.vernier_delay_line_0.stop_strong.n69 VGND 0.11234f
C3734 tdc_0.vernier_delay_line_0.stop_strong.t19 VGND 0.181057f
C3735 tdc_0.vernier_delay_line_0.stop_strong.t5 VGND 0.055955f
C3736 tdc_0.vernier_delay_line_0.stop_strong.n70 VGND 0.413796f
C3737 tdc_0.vernier_delay_line_0.stop_strong.n71 VGND 0.11234f
C3738 tdc_0.vernier_delay_line_0.stop_strong.t29 VGND 0.181057f
C3739 tdc_0.vernier_delay_line_0.stop_strong.t15 VGND 0.055955f
C3740 tdc_0.vernier_delay_line_0.stop_strong.n72 VGND 0.413796f
C3741 tdc_0.vernier_delay_line_0.stop_strong.n73 VGND 0.11234f
C3742 tdc_0.vernier_delay_line_0.stop_strong.t22 VGND 0.181057f
C3743 tdc_0.vernier_delay_line_0.stop_strong.t8 VGND 0.055955f
C3744 tdc_0.vernier_delay_line_0.stop_strong.n74 VGND 0.413796f
C3745 tdc_0.vernier_delay_line_0.stop_strong.n75 VGND 0.11234f
C3746 tdc_0.vernier_delay_line_0.stop_strong.t24 VGND 0.181057f
C3747 tdc_0.vernier_delay_line_0.stop_strong.t10 VGND 0.055955f
C3748 tdc_0.vernier_delay_line_0.stop_strong.n76 VGND 0.413796f
C3749 tdc_0.vernier_delay_line_0.stop_strong.n77 VGND 0.11234f
C3750 tdc_0.vernier_delay_line_0.stop_strong.t18 VGND 0.181057f
C3751 tdc_0.vernier_delay_line_0.stop_strong.t4 VGND 0.055955f
C3752 tdc_0.vernier_delay_line_0.stop_strong.n78 VGND 0.413796f
C3753 tdc_0.vernier_delay_line_0.stop_strong.n79 VGND 0.11234f
C3754 tdc_0.vernier_delay_line_0.stop_strong.t28 VGND 0.181057f
C3755 tdc_0.vernier_delay_line_0.stop_strong.t14 VGND 0.055955f
C3756 tdc_0.vernier_delay_line_0.stop_strong.n80 VGND 0.413796f
C3757 tdc_0.vernier_delay_line_0.stop_strong.n81 VGND 0.11234f
C3758 tdc_0.vernier_delay_line_0.stop_strong.t21 VGND 0.181057f
C3759 tdc_0.vernier_delay_line_0.stop_strong.t7 VGND 0.055955f
C3760 tdc_0.vernier_delay_line_0.stop_strong.n82 VGND 0.413796f
C3761 tdc_0.vernier_delay_line_0.stop_strong.n83 VGND 0.110532f
C3762 tdc_0.vernier_delay_line_0.stop_strong.n84 VGND 1.2768f
C3763 tdc_0.vernier_delay_line_0.stop_strong.t1 VGND 0.055955f
C3764 tdc_0.vernier_delay_line_0.stop_strong.n85 VGND 0.097761f
C3765 tdc_0.vernier_delay_line_0.stop_strong.t31 VGND 0.179153f
C3766 tdc_0.vernier_delay_line_0.stop_strong.n86 VGND 0.326098f
C3767 tdc_0.stop_buffer_0.stop_strong VGND 0.031003f
C3768 a_9330_16954.t4 VGND 0.228995f
C3769 a_9330_16954.t17 VGND 0.093349f
C3770 a_9330_16954.t13 VGND 0.030133f
C3771 a_9330_16954.n0 VGND 0.086421f
C3772 a_9330_16954.t9 VGND 0.093349f
C3773 a_9330_16954.t38 VGND 0.030133f
C3774 a_9330_16954.n1 VGND 0.088816f
C3775 a_9330_16954.t29 VGND 0.093349f
C3776 a_9330_16954.t26 VGND 0.030133f
C3777 a_9330_16954.n2 VGND 0.088354f
C3778 a_9330_16954.n3 VGND 0.389976f
C3779 a_9330_16954.t16 VGND 0.093349f
C3780 a_9330_16954.t12 VGND 0.030133f
C3781 a_9330_16954.n4 VGND 0.088354f
C3782 a_9330_16954.n5 VGND 0.217864f
C3783 a_9330_16954.t35 VGND 0.093349f
C3784 a_9330_16954.t32 VGND 0.030133f
C3785 a_9330_16954.n6 VGND 0.088354f
C3786 a_9330_16954.n7 VGND 0.217864f
C3787 a_9330_16954.t23 VGND 0.093349f
C3788 a_9330_16954.t20 VGND 0.030133f
C3789 a_9330_16954.n8 VGND 0.088354f
C3790 a_9330_16954.n9 VGND 0.217864f
C3791 a_9330_16954.t25 VGND 0.093349f
C3792 a_9330_16954.t22 VGND 0.030133f
C3793 a_9330_16954.n10 VGND 0.088354f
C3794 a_9330_16954.n11 VGND 0.217864f
C3795 a_9330_16954.t11 VGND 0.093349f
C3796 a_9330_16954.t8 VGND 0.030133f
C3797 a_9330_16954.n12 VGND 0.088354f
C3798 a_9330_16954.n13 VGND 0.217864f
C3799 a_9330_16954.t31 VGND 0.093349f
C3800 a_9330_16954.t28 VGND 0.030133f
C3801 a_9330_16954.n14 VGND 0.088354f
C3802 a_9330_16954.n15 VGND 0.217864f
C3803 a_9330_16954.t19 VGND 0.093349f
C3804 a_9330_16954.t15 VGND 0.030133f
C3805 a_9330_16954.n16 VGND 0.088354f
C3806 a_9330_16954.n17 VGND 0.217864f
C3807 a_9330_16954.t37 VGND 0.093349f
C3808 a_9330_16954.t34 VGND 0.030133f
C3809 a_9330_16954.n18 VGND 0.088354f
C3810 a_9330_16954.n19 VGND 0.217864f
C3811 a_9330_16954.t18 VGND 0.093349f
C3812 a_9330_16954.t14 VGND 0.030133f
C3813 a_9330_16954.n20 VGND 0.088354f
C3814 a_9330_16954.n21 VGND 0.217864f
C3815 a_9330_16954.t36 VGND 0.093349f
C3816 a_9330_16954.t33 VGND 0.030133f
C3817 a_9330_16954.n22 VGND 0.088354f
C3818 a_9330_16954.n23 VGND 0.217864f
C3819 a_9330_16954.t24 VGND 0.093349f
C3820 a_9330_16954.t21 VGND 0.030133f
C3821 a_9330_16954.n24 VGND 0.088354f
C3822 a_9330_16954.n25 VGND 0.217864f
C3823 a_9330_16954.t10 VGND 0.093349f
C3824 a_9330_16954.t39 VGND 0.030133f
C3825 a_9330_16954.n26 VGND 0.088354f
C3826 a_9330_16954.n27 VGND 0.217864f
C3827 a_9330_16954.t30 VGND 0.093349f
C3828 a_9330_16954.t27 VGND 0.030133f
C3829 a_9330_16954.n28 VGND 0.088354f
C3830 a_9330_16954.n29 VGND 0.289551f
C3831 a_9330_16954.n30 VGND 0.109352f
C3832 a_9330_16954.n31 VGND 0.42154f
C3833 a_9330_16954.t0 VGND 0.071536f
C3834 a_9330_16954.n32 VGND 0.133321f
C3835 a_9330_16954.t6 VGND 0.231476f
C3836 a_9330_16954.t2 VGND 0.071536f
C3837 a_9330_16954.n33 VGND 0.529025f
C3838 a_9330_16954.n34 VGND 0.22418f
C3839 a_9330_16954.t5 VGND 0.231476f
C3840 a_9330_16954.t1 VGND 0.071536f
C3841 a_9330_16954.n35 VGND 0.538008f
C3842 a_9330_16954.n36 VGND 0.22418f
C3843 a_9330_16954.t3 VGND 0.071536f
C3844 a_9330_16954.n37 VGND 0.529025f
C3845 a_9330_16954.t7 VGND 0.231476f
C3846 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3847 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C3848 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3849 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3850 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.089265f
C3851 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C3852 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3853 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C3854 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.087824f
C3855 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3856 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3857 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.200787f
C3858 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3859 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3860 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3861 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3862 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.107523f
C3863 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3864 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3865 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND 0.019446f
C3866 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 VGND 0.02496f
C3867 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 VGND 0.02496f
C3868 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 VGND 0.074774f
C3869 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VGND 0.048564f
C3870 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VGND 0.154367f
C3871 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 VGND 0.616703f
C3872 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VGND 0.066879f
C3873 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND 0.062029f
C3874 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VGND 0.067105f
C3875 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 VGND 0.065837f
C3876 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 VGND 0.045809f
C3877 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 VGND 0.676981f
C3878 tdc_0.start_buffer_0.start_delay.t8 VGND 0.069408f
C3879 tdc_0.start_buffer_0.start_delay.t15 VGND 0.022142f
C3880 tdc_0.start_buffer_0.start_delay.n0 VGND 0.04868f
C3881 tdc_0.start_buffer_0.start_delay.t14 VGND 0.069408f
C3882 tdc_0.start_buffer_0.start_delay.t12 VGND 0.022142f
C3883 tdc_0.start_buffer_0.start_delay.n1 VGND 0.048366f
C3884 tdc_0.start_buffer_0.start_delay.n2 VGND 0.015598f
C3885 tdc_0.start_buffer_0.start_delay.t13 VGND 0.069408f
C3886 tdc_0.start_buffer_0.start_delay.t11 VGND 0.022142f
C3887 tdc_0.start_buffer_0.start_delay.n3 VGND 0.04868f
C3888 tdc_0.start_buffer_0.start_delay.t10 VGND 0.069408f
C3889 tdc_0.start_buffer_0.start_delay.t9 VGND 0.022142f
C3890 tdc_0.start_buffer_0.start_delay.n4 VGND 0.048366f
C3891 tdc_0.start_buffer_0.start_delay.n5 VGND 0.015431f
C3892 tdc_0.start_buffer_0.start_delay.n6 VGND 0.181697f
C3893 tdc_0.start_buffer_0.start_delay.t6 VGND 0.1725f
C3894 tdc_0.start_buffer_0.start_delay.t2 VGND 0.05331f
C3895 tdc_0.start_buffer_0.start_delay.n7 VGND 0.471528f
C3896 tdc_0.start_buffer_0.start_delay.t7 VGND 0.1725f
C3897 tdc_0.start_buffer_0.start_delay.t3 VGND 0.05331f
C3898 tdc_0.start_buffer_0.start_delay.n8 VGND 0.400932f
C3899 tdc_0.start_buffer_0.start_delay.t5 VGND 0.1725f
C3900 tdc_0.start_buffer_0.start_delay.t1 VGND 0.05331f
C3901 tdc_0.start_buffer_0.start_delay.n9 VGND 0.394238f
C3902 tdc_0.start_buffer_0.start_delay.n10 VGND 0.167063f
C3903 tdc_0.start_buffer_0.start_delay.t4 VGND 0.170686f
C3904 tdc_0.start_buffer_0.start_delay.n11 VGND 0.310685f
C3905 tdc_0.start_buffer_0.start_delay.t0 VGND 0.05331f
C3906 tdc_0.start_buffer_0.start_delay.n12 VGND 0.09314f
C3907 tdc_0.start_buffer_0.start_delay.n13 VGND 0.131763f
C3908 tdc_0.start_buffer_0.start_delay.n14 VGND 0.129117f
C3909 tdc_0.start_buffer_0.start_buff.t15 VGND 0.079205f
C3910 tdc_0.start_buffer_0.start_buff.t12 VGND 0.025267f
C3911 tdc_0.start_buffer_0.start_buff.n0 VGND 0.055193f
C3912 tdc_0.start_buffer_0.start_buff.t11 VGND 0.079205f
C3913 tdc_0.start_buffer_0.start_buff.t20 VGND 0.025267f
C3914 tdc_0.start_buffer_0.start_buff.n1 VGND 0.055551f
C3915 tdc_0.start_buffer_0.start_buff.n2 VGND 0.017803f
C3916 tdc_0.start_buffer_0.start_buff.t19 VGND 0.079205f
C3917 tdc_0.start_buffer_0.start_buff.t17 VGND 0.025267f
C3918 tdc_0.start_buffer_0.start_buff.n3 VGND 0.055551f
C3919 tdc_0.start_buffer_0.start_buff.t13 VGND 0.079205f
C3920 tdc_0.start_buffer_0.start_buff.t23 VGND 0.025267f
C3921 tdc_0.start_buffer_0.start_buff.n4 VGND 0.055193f
C3922 tdc_0.start_buffer_0.start_buff.n5 VGND 0.017609f
C3923 tdc_0.start_buffer_0.start_buff.n6 VGND 0.464807f
C3924 tdc_0.start_buffer_0.start_buff.t9 VGND 0.063388f
C3925 tdc_0.start_buffer_0.start_buff.t8 VGND 0.19187f
C3926 tdc_0.start_buffer_0.start_buff.n7 VGND 0.486972f
C3927 tdc_0.start_buffer_0.start_buff.n8 VGND 0.25373f
C3928 tdc_0.start_buffer_0.start_buff.t5 VGND 0.19187f
C3929 tdc_0.start_buffer_0.start_buff.n9 VGND 0.435589f
C3930 tdc_0.start_buffer_0.start_buff.t10 VGND 0.079384f
C3931 tdc_0.start_buffer_0.start_buff.t22 VGND 0.025625f
C3932 tdc_0.start_buffer_0.start_buff.n10 VGND 0.073493f
C3933 tdc_0.start_buffer_0.start_buff.t21 VGND 0.079384f
C3934 tdc_0.start_buffer_0.start_buff.t18 VGND 0.025625f
C3935 tdc_0.start_buffer_0.start_buff.n11 VGND 0.07553f
C3936 tdc_0.start_buffer_0.start_buff.t16 VGND 0.079384f
C3937 tdc_0.start_buffer_0.start_buff.t14 VGND 0.025625f
C3938 tdc_0.start_buffer_0.start_buff.n12 VGND 0.075137f
C3939 tdc_0.start_buffer_0.start_buff.n13 VGND 0.3926f
C3940 tdc_0.start_buffer_0.start_buff.n14 VGND 0.092517f
C3941 tdc_0.start_buffer_0.start_buff.n15 VGND 0.090637f
C3942 tdc_0.start_buffer_0.start_buff.t1 VGND 0.060835f
C3943 tdc_0.start_buffer_0.start_buff.n16 VGND 0.10659f
C3944 tdc_0.start_buffer_0.start_buff.t6 VGND 0.196849f
C3945 tdc_0.start_buffer_0.start_buff.t2 VGND 0.060835f
C3946 tdc_0.start_buffer_0.start_buff.n17 VGND 0.457525f
C3947 tdc_0.start_buffer_0.start_buff.t4 VGND 0.196849f
C3948 tdc_0.start_buffer_0.start_buff.t0 VGND 0.060835f
C3949 tdc_0.start_buffer_0.start_buff.n18 VGND 0.449886f
C3950 tdc_0.start_buffer_0.start_buff.n19 VGND 0.190644f
C3951 tdc_0.start_buffer_0.start_buff.t7 VGND 0.196849f
C3952 tdc_0.start_buffer_0.start_buff.t3 VGND 0.060835f
C3953 tdc_0.start_buffer_0.start_buff.n20 VGND 0.449886f
C3954 tdc_0.start_buffer_0.start_buff.n21 VGND 0.114821f
C3955 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VGND 0.09757f
C3956 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VGND 0.030153f
C3957 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 VGND 0.265657f
C3958 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 VGND 0.039259f
C3959 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VGND 0.012524f
C3960 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 VGND 0.027534f
C3961 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 VGND 0.039259f
C3962 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 VGND 0.012524f
C3963 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 VGND 0.027357f
C3964 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 VGND 0.008823f
C3965 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VGND 0.039259f
C3966 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 VGND 0.012524f
C3967 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 VGND 0.027534f
C3968 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 VGND 0.039259f
C3969 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 VGND 0.012524f
C3970 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 VGND 0.027357f
C3971 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 VGND 0.008728f
C3972 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 VGND 0.135162f
C3973 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 VGND 0.046129f
C3974 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 VGND 0.046129f
C3975 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 VGND 0.054044f
C3976 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 VGND 0.046129f
C3977 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 VGND 0.046129f
C3978 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 VGND 0.0538f
C3979 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 VGND 0.495704f
C3980 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 VGND 0.119944f
C3981 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 VGND 0.025758f
C3982 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 VGND 0.025758f
C3983 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 VGND 0.055083f
C3984 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 VGND 0.008586f
C3985 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 VGND 0.008586f
C3986 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 VGND 0.01864f
C3987 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 VGND 0.221512f
C3988 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 VGND 0.09757f
C3989 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 VGND 0.030153f
C3990 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 VGND 0.234486f
C3991 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 VGND 0.050613f
C3992 VDPWR.n0 VGND 0.078815f
C3993 VDPWR.t27 VGND 0.050969f
C3994 VDPWR.n1 VGND 0.115444f
C3995 VDPWR.n2 VGND 0.110601f
C3996 VDPWR.n3 VGND 0.110601f
C3997 VDPWR.t472 VGND 0.599415f
C3998 VDPWR.t26 VGND 0.015736f
C3999 VDPWR.n4 VGND 0.095911f
C4000 VDPWR.n5 VGND 0.075149f
C4001 VDPWR.n6 VGND 0.078803f
C4002 VDPWR.t573 VGND 0.050969f
C4003 VDPWR.n7 VGND 0.115444f
C4004 VDPWR.n8 VGND 0.110601f
C4005 VDPWR.n9 VGND 0.110601f
C4006 VDPWR.t77 VGND 0.596797f
C4007 VDPWR.t572 VGND 0.015668f
C4008 VDPWR.n10 VGND 0.095911f
C4009 VDPWR.n11 VGND 0.075149f
C4010 VDPWR.n12 VGND 0.047195f
C4011 VDPWR.t443 VGND 0.05099f
C4012 VDPWR.n13 VGND 0.052839f
C4013 VDPWR.n14 VGND 0.047195f
C4014 VDPWR.n15 VGND 0.03114f
C4015 VDPWR.n16 VGND 0.03114f
C4016 VDPWR.t442 VGND 0.464946f
C4017 VDPWR.n17 VGND 0.25485f
C4018 VDPWR.n18 VGND 0.03114f
C4019 VDPWR.n19 VGND 0.03114f
C4020 VDPWR.n20 VGND 0.047195f
C4021 VDPWR.n21 VGND 0.047195f
C4022 VDPWR.n22 VGND 0.057877f
C4023 VDPWR.t373 VGND 0.013587f
C4024 VDPWR.t23 VGND 0.013587f
C4025 VDPWR.n23 VGND 0.039656f
C4026 VDPWR.t100 VGND 0.050166f
C4027 VDPWR.n24 VGND 0.180877f
C4028 VDPWR.n25 VGND 0.078203f
C4029 VDPWR.n26 VGND 0.057877f
C4030 VDPWR.n27 VGND 0.036626f
C4031 VDPWR.n28 VGND 0.199745f
C4032 VDPWR.t511 VGND 0.170658f
C4033 VDPWR.n29 VGND 0.09447f
C4034 VDPWR.n30 VGND 0.078203f
C4035 VDPWR.t439 VGND 0.097099f
C4036 VDPWR.n31 VGND 0.064732f
C4037 VDPWR.t463 VGND 0.097099f
C4038 VDPWR.t451 VGND 0.191438f
C4039 VDPWR.n32 VGND 0.199745f
C4040 VDPWR.n33 VGND 0.057877f
C4041 VDPWR.t464 VGND 0.013587f
C4042 VDPWR.t440 VGND 0.013587f
C4043 VDPWR.n34 VGND 0.039656f
C4044 VDPWR.t452 VGND 0.050166f
C4045 VDPWR.n35 VGND 0.180877f
C4046 VDPWR.n36 VGND 0.047195f
C4047 VDPWR.t455 VGND 0.05099f
C4048 VDPWR.n37 VGND 0.052839f
C4049 VDPWR.n38 VGND 0.047195f
C4050 VDPWR.n39 VGND 0.03114f
C4051 VDPWR.n40 VGND 0.03114f
C4052 VDPWR.t454 VGND 0.464946f
C4053 VDPWR.n41 VGND 0.25485f
C4054 VDPWR.n42 VGND 0.03114f
C4055 VDPWR.n43 VGND 0.03114f
C4056 VDPWR.n44 VGND 0.049252f
C4057 VDPWR.n45 VGND 0.047195f
C4058 VDPWR.n46 VGND 0.057877f
C4059 VDPWR.t504 VGND 0.013587f
C4060 VDPWR.t502 VGND 0.013587f
C4061 VDPWR.n47 VGND 0.039082f
C4062 VDPWR.t583 VGND 0.050166f
C4063 VDPWR.n48 VGND 0.171056f
C4064 VDPWR.n49 VGND 0.078203f
C4065 VDPWR.n50 VGND 0.057877f
C4066 VDPWR.n51 VGND 0.036626f
C4067 VDPWR.n52 VGND 0.199745f
C4068 VDPWR.t113 VGND 0.170658f
C4069 VDPWR.n53 VGND 0.09447f
C4070 VDPWR.n54 VGND 0.078203f
C4071 VDPWR.t445 VGND 0.097099f
C4072 VDPWR.n55 VGND 0.064732f
C4073 VDPWR.t433 VGND 0.097099f
C4074 VDPWR.t460 VGND 0.191438f
C4075 VDPWR.n56 VGND 0.199745f
C4076 VDPWR.n57 VGND 0.058012f
C4077 VDPWR.t434 VGND 0.013587f
C4078 VDPWR.t446 VGND 0.013587f
C4079 VDPWR.n58 VGND 0.039656f
C4080 VDPWR.t461 VGND 0.050166f
C4081 VDPWR.n59 VGND 0.180877f
C4082 VDPWR.n60 VGND 0.036408f
C4083 VDPWR.n61 VGND 0.033884f
C4084 VDPWR.n62 VGND 0.09447f
C4085 VDPWR.n63 VGND 0.057877f
C4086 VDPWR.n64 VGND 0.036626f
C4087 VDPWR.n65 VGND 0.348672f
C4088 VDPWR.n66 VGND 0.348672f
C4089 VDPWR.t138 VGND 0.170658f
C4090 VDPWR.t503 VGND 0.097099f
C4091 VDPWR.t582 VGND 0.191438f
C4092 VDPWR.t501 VGND 0.097099f
C4093 VDPWR.n67 VGND 0.064732f
C4094 VDPWR.n68 VGND 0.09447f
C4095 VDPWR.n69 VGND 0.09447f
C4096 VDPWR.n70 VGND 0.033884f
C4097 VDPWR.n71 VGND 0.036783f
C4098 VDPWR.n72 VGND 0.044244f
C4099 VDPWR.n73 VGND 0.076499f
C4100 VDPWR.t598 VGND 0.05099f
C4101 VDPWR.n74 VGND 0.04954f
C4102 VDPWR.n75 VGND 0.094073f
C4103 VDPWR.n76 VGND 0.012369f
C4104 VDPWR.n77 VGND 0.061487f
C4105 VDPWR.n78 VGND 0.061487f
C4106 VDPWR.n79 VGND 0.344359f
C4107 VDPWR.n80 VGND 0.061487f
C4108 VDPWR.n81 VGND 0.061487f
C4109 VDPWR.n82 VGND 0.014168f
C4110 VDPWR.n83 VGND 0.094073f
C4111 VDPWR.n84 VGND 0.054612f
C4112 VDPWR.t453 VGND 0.020756f
C4113 VDPWR.t616 VGND 0.0067f
C4114 VDPWR.n85 VGND 0.020461f
C4115 VDPWR.t432 VGND 0.020475f
C4116 VDPWR.t459 VGND 0.022151f
C4117 VDPWR.n86 VGND 0.021732f
C4118 VDPWR.t444 VGND 0.022076f
C4119 VDPWR.n87 VGND 0.015124f
C4120 VDPWR.t618 VGND 0.006419f
C4121 VDPWR.t619 VGND 0.008239f
C4122 VDPWR.t627 VGND 0.008239f
C4123 VDPWR.n88 VGND 0.024694f
C4124 VDPWR.n89 VGND 0.15186f
C4125 VDPWR.n90 VGND 0.122334f
C4126 VDPWR.n91 VGND 0.149158f
C4127 VDPWR.n92 VGND 0.042752f
C4128 VDPWR.n93 VGND 0.037122f
C4129 VDPWR.n94 VGND 0.036408f
C4130 VDPWR.n95 VGND 0.033884f
C4131 VDPWR.n96 VGND 0.09447f
C4132 VDPWR.n97 VGND 0.057877f
C4133 VDPWR.n98 VGND 0.036626f
C4134 VDPWR.n99 VGND 0.348672f
C4135 VDPWR.n100 VGND 0.348672f
C4136 VDPWR.t102 VGND 0.170658f
C4137 VDPWR.t372 VGND 0.097099f
C4138 VDPWR.t99 VGND 0.191438f
C4139 VDPWR.t22 VGND 0.097099f
C4140 VDPWR.n101 VGND 0.064732f
C4141 VDPWR.n102 VGND 0.09447f
C4142 VDPWR.n103 VGND 0.09447f
C4143 VDPWR.n104 VGND 0.033884f
C4144 VDPWR.n105 VGND 0.036783f
C4145 VDPWR.n106 VGND 0.044244f
C4146 VDPWR.n107 VGND 0.074573f
C4147 VDPWR.t485 VGND 0.05099f
C4148 VDPWR.n108 VGND 0.04954f
C4149 VDPWR.n109 VGND 0.094073f
C4150 VDPWR.n110 VGND 0.014168f
C4151 VDPWR.n111 VGND 0.061487f
C4152 VDPWR.n112 VGND 0.061487f
C4153 VDPWR.n113 VGND 0.344359f
C4154 VDPWR.n114 VGND 0.061487f
C4155 VDPWR.n115 VGND 0.061487f
C4156 VDPWR.n116 VGND 0.014168f
C4157 VDPWR.n117 VGND 0.094073f
C4158 VDPWR.n118 VGND 0.055663f
C4159 VDPWR.t441 VGND 0.020756f
C4160 VDPWR.t620 VGND 0.0067f
C4161 VDPWR.n119 VGND 0.020472f
C4162 VDPWR.t462 VGND 0.020475f
C4163 VDPWR.t450 VGND 0.022151f
C4164 VDPWR.n120 VGND 0.021732f
C4165 VDPWR.t438 VGND 0.022076f
C4166 VDPWR.n121 VGND 0.015124f
C4167 VDPWR.t622 VGND 0.006419f
C4168 VDPWR.t625 VGND 0.008239f
C4169 VDPWR.t628 VGND 0.008239f
C4170 VDPWR.n122 VGND 0.024694f
C4171 VDPWR.n123 VGND 0.15186f
C4172 VDPWR.n124 VGND 0.121787f
C4173 VDPWR.n125 VGND 0.149694f
C4174 VDPWR.n126 VGND 0.029594f
C4175 VDPWR.n127 VGND 0.030252f
C4176 VDPWR.t78 VGND 0.050974f
C4177 VDPWR.n128 VGND 0.119109f
C4178 VDPWR.n129 VGND 0.239269f
C4179 VDPWR.n130 VGND 0.058006f
C4180 VDPWR.n131 VGND 0.041651f
C4181 VDPWR.n132 VGND 0.311313f
C4182 VDPWR.n133 VGND 0.025446f
C4183 VDPWR.n134 VGND 0.535617f
C4184 VDPWR.n135 VGND 0.100578f
C4185 VDPWR.n136 VGND 0.024738f
C4186 VDPWR.n137 VGND 0.110649f
C4187 VDPWR.n138 VGND 0.072182f
C4188 VDPWR.t473 VGND 0.050974f
C4189 VDPWR.n139 VGND 0.119109f
C4190 VDPWR.n140 VGND 0.117419f
C4191 VDPWR.n141 VGND 0.058006f
C4192 VDPWR.n142 VGND 0.041651f
C4193 VDPWR.n143 VGND 0.312713f
C4194 VDPWR.n144 VGND 0.025434f
C4195 VDPWR.n145 VGND 0.537491f
C4196 VDPWR.n146 VGND 0.100578f
C4197 VDPWR.n147 VGND 0.024738f
C4198 VDPWR.n148 VGND 0.110649f
C4199 VDPWR.n149 VGND 0.072182f
C4200 VDPWR.n150 VGND 0.107712f
C4201 VDPWR.n151 VGND 0.051562f
C4202 VDPWR.t332 VGND 0.05099f
C4203 VDPWR.n152 VGND 0.140617f
C4204 VDPWR.n153 VGND 0.225436f
C4205 VDPWR.t331 VGND 0.232473f
C4206 VDPWR.n154 VGND 0.03114f
C4207 VDPWR.n155 VGND 0.135655f
C4208 VDPWR.n156 VGND 0.019839f
C4209 VDPWR.n157 VGND 0.061493f
C4210 VDPWR.n158 VGND 0.061487f
C4211 VDPWR.n159 VGND 0.003523f
C4212 VDPWR.n160 VGND 0.073016f
C4213 VDPWR.n161 VGND 0.101812f
C4214 VDPWR.t534 VGND 0.051124f
C4215 VDPWR.n162 VGND 0.099892f
C4216 VDPWR.n163 VGND 0.076349f
C4217 VDPWR.n164 VGND 0.30266f
C4218 VDPWR.t139 VGND 0.285828f
C4219 VDPWR.t140 VGND 0.051124f
C4220 VDPWR.n165 VGND 0.010355f
C4221 VDPWR.n166 VGND 0.099892f
C4222 VDPWR.t621 VGND 0.015661f
C4223 VDPWR.t624 VGND 0.021113f
C4224 VDPWR.n167 VGND 0.023494f
C4225 VDPWR.n168 VGND 0.100362f
C4226 VDPWR.n169 VGND 0.078815f
C4227 VDPWR.t1 VGND 0.050969f
C4228 VDPWR.n170 VGND 0.115444f
C4229 VDPWR.n171 VGND 0.110601f
C4230 VDPWR.n172 VGND 0.110601f
C4231 VDPWR.t178 VGND 0.599415f
C4232 VDPWR.t0 VGND 0.015736f
C4233 VDPWR.n173 VGND 0.095911f
C4234 VDPWR.n174 VGND 0.075149f
C4235 VDPWR.n175 VGND 0.078803f
C4236 VDPWR.t21 VGND 0.050969f
C4237 VDPWR.n176 VGND 0.115444f
C4238 VDPWR.n177 VGND 0.110601f
C4239 VDPWR.n178 VGND 0.110601f
C4240 VDPWR.t222 VGND 0.596797f
C4241 VDPWR.t20 VGND 0.015668f
C4242 VDPWR.n179 VGND 0.095911f
C4243 VDPWR.n180 VGND 0.075149f
C4244 VDPWR.n181 VGND 0.047195f
C4245 VDPWR.t340 VGND 0.05099f
C4246 VDPWR.n182 VGND 0.052839f
C4247 VDPWR.n183 VGND 0.047195f
C4248 VDPWR.n184 VGND 0.03114f
C4249 VDPWR.n185 VGND 0.03114f
C4250 VDPWR.t339 VGND 0.464946f
C4251 VDPWR.n186 VGND 0.25485f
C4252 VDPWR.n187 VGND 0.03114f
C4253 VDPWR.n188 VGND 0.03114f
C4254 VDPWR.n189 VGND 0.047195f
C4255 VDPWR.n190 VGND 0.047195f
C4256 VDPWR.n191 VGND 0.057877f
C4257 VDPWR.t328 VGND 0.013587f
C4258 VDPWR.t562 VGND 0.013587f
C4259 VDPWR.n192 VGND 0.039656f
C4260 VDPWR.t560 VGND 0.050166f
C4261 VDPWR.n193 VGND 0.180877f
C4262 VDPWR.n194 VGND 0.078203f
C4263 VDPWR.n195 VGND 0.057877f
C4264 VDPWR.n196 VGND 0.036626f
C4265 VDPWR.n197 VGND 0.199745f
C4266 VDPWR.t199 VGND 0.170658f
C4267 VDPWR.n198 VGND 0.09447f
C4268 VDPWR.n199 VGND 0.078203f
C4269 VDPWR.t418 VGND 0.097099f
C4270 VDPWR.n200 VGND 0.064732f
C4271 VDPWR.t354 VGND 0.097099f
C4272 VDPWR.t196 VGND 0.191438f
C4273 VDPWR.n201 VGND 0.199745f
C4274 VDPWR.n202 VGND 0.057877f
C4275 VDPWR.t355 VGND 0.013587f
C4276 VDPWR.t419 VGND 0.013587f
C4277 VDPWR.n203 VGND 0.039656f
C4278 VDPWR.t197 VGND 0.050166f
C4279 VDPWR.n204 VGND 0.180877f
C4280 VDPWR.n205 VGND 0.047195f
C4281 VDPWR.t137 VGND 0.05099f
C4282 VDPWR.n206 VGND 0.052839f
C4283 VDPWR.n207 VGND 0.047195f
C4284 VDPWR.n208 VGND 0.03114f
C4285 VDPWR.n209 VGND 0.03114f
C4286 VDPWR.t136 VGND 0.464946f
C4287 VDPWR.n210 VGND 0.25485f
C4288 VDPWR.n211 VGND 0.03114f
C4289 VDPWR.n212 VGND 0.03114f
C4290 VDPWR.n213 VGND 0.047195f
C4291 VDPWR.n214 VGND 0.047195f
C4292 VDPWR.n215 VGND 0.057877f
C4293 VDPWR.t508 VGND 0.013587f
C4294 VDPWR.t131 VGND 0.013587f
C4295 VDPWR.n216 VGND 0.039656f
C4296 VDPWR.t427 VGND 0.050166f
C4297 VDPWR.n217 VGND 0.180877f
C4298 VDPWR.n218 VGND 0.078203f
C4299 VDPWR.n219 VGND 0.057877f
C4300 VDPWR.n220 VGND 0.036626f
C4301 VDPWR.n221 VGND 0.199745f
C4302 VDPWR.t509 VGND 0.170658f
C4303 VDPWR.n222 VGND 0.09447f
C4304 VDPWR.n223 VGND 0.078203f
C4305 VDPWR.t134 VGND 0.097099f
C4306 VDPWR.n224 VGND 0.064732f
C4307 VDPWR.t165 VGND 0.097099f
C4308 VDPWR.t163 VGND 0.191438f
C4309 VDPWR.n225 VGND 0.199745f
C4310 VDPWR.n226 VGND 0.057877f
C4311 VDPWR.t166 VGND 0.013587f
C4312 VDPWR.t135 VGND 0.013587f
C4313 VDPWR.n227 VGND 0.039656f
C4314 VDPWR.t164 VGND 0.050166f
C4315 VDPWR.n228 VGND 0.180877f
C4316 VDPWR.n229 VGND 0.047195f
C4317 VDPWR.t567 VGND 0.05099f
C4318 VDPWR.n230 VGND 0.052839f
C4319 VDPWR.n231 VGND 0.047195f
C4320 VDPWR.n232 VGND 0.03114f
C4321 VDPWR.n233 VGND 0.03114f
C4322 VDPWR.t386 VGND 0.464946f
C4323 VDPWR.n234 VGND 0.25485f
C4324 VDPWR.n235 VGND 0.03114f
C4325 VDPWR.n236 VGND 0.03114f
C4326 VDPWR.n237 VGND 0.047195f
C4327 VDPWR.n238 VGND 0.047195f
C4328 VDPWR.n239 VGND 0.057877f
C4329 VDPWR.t244 VGND 0.013587f
C4330 VDPWR.t242 VGND 0.013587f
C4331 VDPWR.n240 VGND 0.039656f
C4332 VDPWR.t284 VGND 0.050166f
C4333 VDPWR.n241 VGND 0.180877f
C4334 VDPWR.n242 VGND 0.078203f
C4335 VDPWR.n243 VGND 0.057877f
C4336 VDPWR.n244 VGND 0.036626f
C4337 VDPWR.n245 VGND 0.199745f
C4338 VDPWR.t558 VGND 0.170658f
C4339 VDPWR.n246 VGND 0.09447f
C4340 VDPWR.n247 VGND 0.078203f
C4341 VDPWR.t337 VGND 0.097099f
C4342 VDPWR.n248 VGND 0.064732f
C4343 VDPWR.t590 VGND 0.097099f
C4344 VDPWR.t592 VGND 0.191438f
C4345 VDPWR.n249 VGND 0.199745f
C4346 VDPWR.n250 VGND 0.057877f
C4347 VDPWR.t591 VGND 0.013587f
C4348 VDPWR.t338 VGND 0.013587f
C4349 VDPWR.n251 VGND 0.039656f
C4350 VDPWR.t593 VGND 0.050166f
C4351 VDPWR.n252 VGND 0.180877f
C4352 VDPWR.n253 VGND 0.047195f
C4353 VDPWR.t553 VGND 0.05099f
C4354 VDPWR.n254 VGND 0.052839f
C4355 VDPWR.n255 VGND 0.047195f
C4356 VDPWR.n256 VGND 0.03114f
C4357 VDPWR.n257 VGND 0.03114f
C4358 VDPWR.t250 VGND 0.464946f
C4359 VDPWR.n258 VGND 0.25485f
C4360 VDPWR.n259 VGND 0.03114f
C4361 VDPWR.n260 VGND 0.03114f
C4362 VDPWR.n261 VGND 0.047195f
C4363 VDPWR.n262 VGND 0.047195f
C4364 VDPWR.n263 VGND 0.057877f
C4365 VDPWR.t515 VGND 0.013587f
C4366 VDPWR.t336 VGND 0.013587f
C4367 VDPWR.n264 VGND 0.039656f
C4368 VDPWR.t334 VGND 0.050166f
C4369 VDPWR.n265 VGND 0.180877f
C4370 VDPWR.n266 VGND 0.078203f
C4371 VDPWR.n267 VGND 0.057877f
C4372 VDPWR.n268 VGND 0.036626f
C4373 VDPWR.n269 VGND 0.199745f
C4374 VDPWR.t226 VGND 0.170658f
C4375 VDPWR.n270 VGND 0.09447f
C4376 VDPWR.n271 VGND 0.078203f
C4377 VDPWR.t285 VGND 0.097099f
C4378 VDPWR.n272 VGND 0.064732f
C4379 VDPWR.t416 VGND 0.097099f
C4380 VDPWR.t301 VGND 0.191438f
C4381 VDPWR.n273 VGND 0.199745f
C4382 VDPWR.n274 VGND 0.057877f
C4383 VDPWR.t417 VGND 0.013587f
C4384 VDPWR.t286 VGND 0.013587f
C4385 VDPWR.n275 VGND 0.039656f
C4386 VDPWR.t302 VGND 0.050166f
C4387 VDPWR.n276 VGND 0.180877f
C4388 VDPWR.n277 VGND 0.047195f
C4389 VDPWR.t612 VGND 0.05099f
C4390 VDPWR.n278 VGND 0.052839f
C4391 VDPWR.n279 VGND 0.047195f
C4392 VDPWR.n280 VGND 0.03114f
C4393 VDPWR.n281 VGND 0.03114f
C4394 VDPWR.t367 VGND 0.464946f
C4395 VDPWR.n282 VGND 0.25485f
C4396 VDPWR.n283 VGND 0.03114f
C4397 VDPWR.n284 VGND 0.03114f
C4398 VDPWR.n285 VGND 0.047195f
C4399 VDPWR.n286 VGND 0.047195f
C4400 VDPWR.n287 VGND 0.057877f
C4401 VDPWR.t207 VGND 0.013587f
C4402 VDPWR.t221 VGND 0.013587f
C4403 VDPWR.n288 VGND 0.039656f
C4404 VDPWR.t209 VGND 0.050166f
C4405 VDPWR.n289 VGND 0.180877f
C4406 VDPWR.n290 VGND 0.078203f
C4407 VDPWR.n291 VGND 0.057877f
C4408 VDPWR.n292 VGND 0.036626f
C4409 VDPWR.n293 VGND 0.199745f
C4410 VDPWR.t3 VGND 0.170658f
C4411 VDPWR.n294 VGND 0.09447f
C4412 VDPWR.n295 VGND 0.078203f
C4413 VDPWR.t29 VGND 0.097099f
C4414 VDPWR.n296 VGND 0.064732f
C4415 VDPWR.t97 VGND 0.097099f
C4416 VDPWR.t610 VGND 0.191438f
C4417 VDPWR.n297 VGND 0.199745f
C4418 VDPWR.n298 VGND 0.057877f
C4419 VDPWR.t98 VGND 0.013587f
C4420 VDPWR.t30 VGND 0.013587f
C4421 VDPWR.n299 VGND 0.039656f
C4422 VDPWR.t611 VGND 0.050166f
C4423 VDPWR.n300 VGND 0.180877f
C4424 VDPWR.n301 VGND 0.047195f
C4425 VDPWR.t467 VGND 0.05099f
C4426 VDPWR.n302 VGND 0.052839f
C4427 VDPWR.n303 VGND 0.047195f
C4428 VDPWR.n304 VGND 0.03114f
C4429 VDPWR.n305 VGND 0.03114f
C4430 VDPWR.t466 VGND 0.464946f
C4431 VDPWR.n306 VGND 0.25485f
C4432 VDPWR.n307 VGND 0.03114f
C4433 VDPWR.n308 VGND 0.03114f
C4434 VDPWR.n309 VGND 0.047195f
C4435 VDPWR.n310 VGND 0.047195f
C4436 VDPWR.n311 VGND 0.057877f
C4437 VDPWR.t513 VGND 0.013587f
C4438 VDPWR.t149 VGND 0.013587f
C4439 VDPWR.n312 VGND 0.039656f
C4440 VDPWR.t330 VGND 0.050166f
C4441 VDPWR.n313 VGND 0.180877f
C4442 VDPWR.n314 VGND 0.078203f
C4443 VDPWR.n315 VGND 0.057877f
C4444 VDPWR.n316 VGND 0.036626f
C4445 VDPWR.n317 VGND 0.199745f
C4446 VDPWR.t112 VGND 0.170658f
C4447 VDPWR.n318 VGND 0.09447f
C4448 VDPWR.n319 VGND 0.078203f
C4449 VDPWR.t448 VGND 0.097099f
C4450 VDPWR.n320 VGND 0.064732f
C4451 VDPWR.t436 VGND 0.097099f
C4452 VDPWR.t457 VGND 0.191438f
C4453 VDPWR.n321 VGND 0.199745f
C4454 VDPWR.n322 VGND 0.058012f
C4455 VDPWR.t437 VGND 0.013587f
C4456 VDPWR.t449 VGND 0.013587f
C4457 VDPWR.n323 VGND 0.039656f
C4458 VDPWR.t458 VGND 0.050166f
C4459 VDPWR.n324 VGND 0.180877f
C4460 VDPWR.n325 VGND 0.036408f
C4461 VDPWR.n326 VGND 0.033884f
C4462 VDPWR.n327 VGND 0.09447f
C4463 VDPWR.n328 VGND 0.057877f
C4464 VDPWR.n329 VGND 0.036626f
C4465 VDPWR.n330 VGND 0.348672f
C4466 VDPWR.n331 VGND 0.348672f
C4467 VDPWR.t520 VGND 0.170658f
C4468 VDPWR.t512 VGND 0.097099f
C4469 VDPWR.t329 VGND 0.191438f
C4470 VDPWR.t148 VGND 0.097099f
C4471 VDPWR.n332 VGND 0.064732f
C4472 VDPWR.n333 VGND 0.09447f
C4473 VDPWR.n334 VGND 0.09447f
C4474 VDPWR.n335 VGND 0.033884f
C4475 VDPWR.n336 VGND 0.036783f
C4476 VDPWR.n337 VGND 0.044244f
C4477 VDPWR.n338 VGND 0.074573f
C4478 VDPWR.t579 VGND 0.05099f
C4479 VDPWR.n339 VGND 0.04954f
C4480 VDPWR.n340 VGND 0.094073f
C4481 VDPWR.n341 VGND 0.014168f
C4482 VDPWR.n342 VGND 0.061487f
C4483 VDPWR.n343 VGND 0.061487f
C4484 VDPWR.n344 VGND 0.344359f
C4485 VDPWR.n345 VGND 0.061487f
C4486 VDPWR.n346 VGND 0.061487f
C4487 VDPWR.n347 VGND 0.014168f
C4488 VDPWR.n348 VGND 0.094073f
C4489 VDPWR.n349 VGND 0.054288f
C4490 VDPWR.t465 VGND 0.020756f
C4491 VDPWR.t615 VGND 0.0067f
C4492 VDPWR.n350 VGND 0.020458f
C4493 VDPWR.t435 VGND 0.020475f
C4494 VDPWR.t456 VGND 0.022151f
C4495 VDPWR.n351 VGND 0.021732f
C4496 VDPWR.t447 VGND 0.022076f
C4497 VDPWR.n352 VGND 0.015124f
C4498 VDPWR.t626 VGND 0.006419f
C4499 VDPWR.t617 VGND 0.008239f
C4500 VDPWR.t623 VGND 0.008239f
C4501 VDPWR.n353 VGND 0.024694f
C4502 VDPWR.n354 VGND 0.15186f
C4503 VDPWR.n355 VGND 0.122498f
C4504 VDPWR.n356 VGND 0.148997f
C4505 VDPWR.n357 VGND 0.042795f
C4506 VDPWR.n358 VGND 0.037122f
C4507 VDPWR.n359 VGND 0.036408f
C4508 VDPWR.n360 VGND 0.033884f
C4509 VDPWR.n361 VGND 0.09447f
C4510 VDPWR.n362 VGND 0.057877f
C4511 VDPWR.n363 VGND 0.036626f
C4512 VDPWR.n364 VGND 0.348672f
C4513 VDPWR.n365 VGND 0.348672f
C4514 VDPWR.t390 VGND 0.170658f
C4515 VDPWR.t206 VGND 0.097099f
C4516 VDPWR.t208 VGND 0.191438f
C4517 VDPWR.t220 VGND 0.097099f
C4518 VDPWR.n366 VGND 0.064732f
C4519 VDPWR.n367 VGND 0.09447f
C4520 VDPWR.n368 VGND 0.09447f
C4521 VDPWR.n369 VGND 0.033884f
C4522 VDPWR.n370 VGND 0.036783f
C4523 VDPWR.n371 VGND 0.044244f
C4524 VDPWR.n372 VGND 0.074573f
C4525 VDPWR.t368 VGND 0.05099f
C4526 VDPWR.n373 VGND 0.04954f
C4527 VDPWR.n374 VGND 0.094073f
C4528 VDPWR.n375 VGND 0.014168f
C4529 VDPWR.n376 VGND 0.061487f
C4530 VDPWR.n377 VGND 0.061487f
C4531 VDPWR.n378 VGND 0.344359f
C4532 VDPWR.n379 VGND 0.061487f
C4533 VDPWR.n380 VGND 0.061487f
C4534 VDPWR.n381 VGND 0.014168f
C4535 VDPWR.n382 VGND 0.094073f
C4536 VDPWR.n383 VGND 0.083636f
C4537 VDPWR.n384 VGND 0.037122f
C4538 VDPWR.n385 VGND 0.036408f
C4539 VDPWR.n386 VGND 0.033884f
C4540 VDPWR.n387 VGND 0.09447f
C4541 VDPWR.n388 VGND 0.057877f
C4542 VDPWR.n389 VGND 0.036626f
C4543 VDPWR.n390 VGND 0.348672f
C4544 VDPWR.n391 VGND 0.348672f
C4545 VDPWR.t129 VGND 0.170658f
C4546 VDPWR.t514 VGND 0.097099f
C4547 VDPWR.t333 VGND 0.191438f
C4548 VDPWR.t335 VGND 0.097099f
C4549 VDPWR.n392 VGND 0.064732f
C4550 VDPWR.n393 VGND 0.09447f
C4551 VDPWR.n394 VGND 0.09447f
C4552 VDPWR.n395 VGND 0.033884f
C4553 VDPWR.n396 VGND 0.036783f
C4554 VDPWR.n397 VGND 0.044244f
C4555 VDPWR.n398 VGND 0.074573f
C4556 VDPWR.t251 VGND 0.05099f
C4557 VDPWR.n399 VGND 0.04954f
C4558 VDPWR.n400 VGND 0.094073f
C4559 VDPWR.n401 VGND 0.014168f
C4560 VDPWR.n402 VGND 0.061487f
C4561 VDPWR.n403 VGND 0.061487f
C4562 VDPWR.n404 VGND 0.344359f
C4563 VDPWR.n405 VGND 0.061487f
C4564 VDPWR.n406 VGND 0.061487f
C4565 VDPWR.n407 VGND 0.014168f
C4566 VDPWR.n408 VGND 0.094073f
C4567 VDPWR.n409 VGND 0.083636f
C4568 VDPWR.n410 VGND 0.037122f
C4569 VDPWR.n411 VGND 0.036408f
C4570 VDPWR.n412 VGND 0.033884f
C4571 VDPWR.n413 VGND 0.09447f
C4572 VDPWR.n414 VGND 0.057877f
C4573 VDPWR.n415 VGND 0.036626f
C4574 VDPWR.n416 VGND 0.348672f
C4575 VDPWR.n417 VGND 0.348672f
C4576 VDPWR.t171 VGND 0.170658f
C4577 VDPWR.t243 VGND 0.097099f
C4578 VDPWR.t283 VGND 0.191438f
C4579 VDPWR.t241 VGND 0.097099f
C4580 VDPWR.n418 VGND 0.064732f
C4581 VDPWR.n419 VGND 0.09447f
C4582 VDPWR.n420 VGND 0.09447f
C4583 VDPWR.n421 VGND 0.033884f
C4584 VDPWR.n422 VGND 0.036783f
C4585 VDPWR.n423 VGND 0.044244f
C4586 VDPWR.n424 VGND 0.074573f
C4587 VDPWR.t387 VGND 0.05099f
C4588 VDPWR.n425 VGND 0.04954f
C4589 VDPWR.n426 VGND 0.094073f
C4590 VDPWR.n427 VGND 0.014168f
C4591 VDPWR.n428 VGND 0.061487f
C4592 VDPWR.n429 VGND 0.061487f
C4593 VDPWR.n430 VGND 0.344359f
C4594 VDPWR.n431 VGND 0.061487f
C4595 VDPWR.n432 VGND 0.061487f
C4596 VDPWR.n433 VGND 0.014168f
C4597 VDPWR.n434 VGND 0.094073f
C4598 VDPWR.n435 VGND 0.083636f
C4599 VDPWR.n436 VGND 0.037122f
C4600 VDPWR.n437 VGND 0.036408f
C4601 VDPWR.n438 VGND 0.033884f
C4602 VDPWR.n439 VGND 0.09447f
C4603 VDPWR.n440 VGND 0.057877f
C4604 VDPWR.n441 VGND 0.036626f
C4605 VDPWR.n442 VGND 0.348672f
C4606 VDPWR.n443 VGND 0.348672f
C4607 VDPWR.t491 VGND 0.170658f
C4608 VDPWR.t507 VGND 0.097099f
C4609 VDPWR.t426 VGND 0.191438f
C4610 VDPWR.t130 VGND 0.097099f
C4611 VDPWR.n444 VGND 0.064732f
C4612 VDPWR.n445 VGND 0.09447f
C4613 VDPWR.n446 VGND 0.09447f
C4614 VDPWR.n447 VGND 0.033884f
C4615 VDPWR.n448 VGND 0.036783f
C4616 VDPWR.n449 VGND 0.044244f
C4617 VDPWR.n450 VGND 0.074573f
C4618 VDPWR.t605 VGND 0.05099f
C4619 VDPWR.n451 VGND 0.04954f
C4620 VDPWR.n452 VGND 0.094073f
C4621 VDPWR.n453 VGND 0.014168f
C4622 VDPWR.n454 VGND 0.061487f
C4623 VDPWR.n455 VGND 0.061487f
C4624 VDPWR.n456 VGND 0.344359f
C4625 VDPWR.n457 VGND 0.061487f
C4626 VDPWR.n458 VGND 0.061487f
C4627 VDPWR.n459 VGND 0.014168f
C4628 VDPWR.n460 VGND 0.094073f
C4629 VDPWR.n461 VGND 0.083636f
C4630 VDPWR.n462 VGND 0.037122f
C4631 VDPWR.n463 VGND 0.036408f
C4632 VDPWR.n464 VGND 0.033884f
C4633 VDPWR.n465 VGND 0.09447f
C4634 VDPWR.n466 VGND 0.057877f
C4635 VDPWR.n467 VGND 0.036626f
C4636 VDPWR.n468 VGND 0.348672f
C4637 VDPWR.n469 VGND 0.348672f
C4638 VDPWR.t606 VGND 0.170658f
C4639 VDPWR.t327 VGND 0.097099f
C4640 VDPWR.t559 VGND 0.191438f
C4641 VDPWR.t561 VGND 0.097099f
C4642 VDPWR.n470 VGND 0.064732f
C4643 VDPWR.n471 VGND 0.09447f
C4644 VDPWR.n472 VGND 0.09447f
C4645 VDPWR.n473 VGND 0.033884f
C4646 VDPWR.n474 VGND 0.036783f
C4647 VDPWR.n475 VGND 0.044244f
C4648 VDPWR.n476 VGND 0.074573f
C4649 VDPWR.t589 VGND 0.05099f
C4650 VDPWR.n477 VGND 0.04954f
C4651 VDPWR.n478 VGND 0.094073f
C4652 VDPWR.n479 VGND 0.014168f
C4653 VDPWR.n480 VGND 0.061487f
C4654 VDPWR.n481 VGND 0.061487f
C4655 VDPWR.n482 VGND 0.344359f
C4656 VDPWR.n483 VGND 0.061487f
C4657 VDPWR.n484 VGND 0.061487f
C4658 VDPWR.n485 VGND 0.014168f
C4659 VDPWR.n486 VGND 0.094073f
C4660 VDPWR.n487 VGND 0.068603f
C4661 VDPWR.n488 VGND 0.046531f
C4662 VDPWR.t223 VGND 0.050974f
C4663 VDPWR.n489 VGND 0.119109f
C4664 VDPWR.n490 VGND 0.221568f
C4665 VDPWR.n491 VGND 0.058006f
C4666 VDPWR.n492 VGND 0.041651f
C4667 VDPWR.n493 VGND 0.311313f
C4668 VDPWR.n494 VGND 0.025446f
C4669 VDPWR.n495 VGND 0.535617f
C4670 VDPWR.n496 VGND 0.100578f
C4671 VDPWR.n497 VGND 0.024738f
C4672 VDPWR.n498 VGND 0.110649f
C4673 VDPWR.n499 VGND 0.072182f
C4674 VDPWR.t179 VGND 0.050974f
C4675 VDPWR.n500 VGND 0.119109f
C4676 VDPWR.n501 VGND 0.117419f
C4677 VDPWR.n502 VGND 0.058006f
C4678 VDPWR.n503 VGND 0.041651f
C4679 VDPWR.n504 VGND 0.312713f
C4680 VDPWR.n505 VGND 0.025434f
C4681 VDPWR.n506 VGND 0.537491f
C4682 VDPWR.n507 VGND 0.100578f
C4683 VDPWR.n508 VGND 0.024738f
C4684 VDPWR.n509 VGND 0.110649f
C4685 VDPWR.n510 VGND 0.072182f
C4686 VDPWR.n511 VGND 1.09207f
C4687 VDPWR.t401 VGND 0.051359f
C4688 VDPWR.t347 VGND 0.050988f
C4689 VDPWR.n512 VGND 0.189533f
C4690 VDPWR.t72 VGND 0.050988f
C4691 VDPWR.n513 VGND 0.100448f
C4692 VDPWR.t490 VGND 0.050988f
C4693 VDPWR.n514 VGND 0.095922f
C4694 VDPWR.n515 VGND 0.062776f
C4695 VDPWR.n516 VGND 0.037653f
C4696 VDPWR.t258 VGND 0.051359f
C4697 VDPWR.t219 VGND 0.050988f
C4698 VDPWR.n517 VGND 0.189533f
C4699 VDPWR.t478 VGND 0.050988f
C4700 VDPWR.n518 VGND 0.100448f
C4701 VDPWR.t215 VGND 0.050988f
C4702 VDPWR.n519 VGND 0.095922f
C4703 VDPWR.n520 VGND 0.062776f
C4704 VDPWR.n521 VGND 0.037653f
C4705 VDPWR.t488 VGND 0.051359f
C4706 VDPWR.t316 VGND 0.050988f
C4707 VDPWR.n522 VGND 0.189533f
C4708 VDPWR.t321 VGND 0.050988f
C4709 VDPWR.n523 VGND 0.100448f
C4710 VDPWR.t378 VGND 0.050988f
C4711 VDPWR.n524 VGND 0.095922f
C4712 VDPWR.n525 VGND 0.062776f
C4713 VDPWR.n526 VGND 0.037653f
C4714 VDPWR.t259 VGND 0.051359f
C4715 VDPWR.t187 VGND 0.050988f
C4716 VDPWR.n527 VGND 0.189533f
C4717 VDPWR.t360 VGND 0.050988f
C4718 VDPWR.n528 VGND 0.100448f
C4719 VDPWR.t489 VGND 0.050988f
C4720 VDPWR.n529 VGND 0.095922f
C4721 VDPWR.n530 VGND 0.062776f
C4722 VDPWR.n531 VGND 0.037653f
C4723 VDPWR.t124 VGND 0.051359f
C4724 VDPWR.t144 VGND 0.050988f
C4725 VDPWR.n532 VGND 0.189533f
C4726 VDPWR.t123 VGND 0.050988f
C4727 VDPWR.n533 VGND 0.100448f
C4728 VDPWR.t216 VGND 0.050988f
C4729 VDPWR.n534 VGND 0.095922f
C4730 VDPWR.n535 VGND 0.062776f
C4731 VDPWR.n536 VGND 0.037653f
C4732 VDPWR.t525 VGND 0.051359f
C4733 VDPWR.t479 VGND 0.050988f
C4734 VDPWR.n537 VGND 0.189533f
C4735 VDPWR.t247 VGND 0.050988f
C4736 VDPWR.n538 VGND 0.100448f
C4737 VDPWR.t492 VGND 0.050988f
C4738 VDPWR.n539 VGND 0.095922f
C4739 VDPWR.n540 VGND 0.062776f
C4740 VDPWR.n541 VGND 0.037653f
C4741 VDPWR.t532 VGND 0.051359f
C4742 VDPWR.t261 VGND 0.050988f
C4743 VDPWR.n542 VGND 0.189533f
C4744 VDPWR.t371 VGND 0.050988f
C4745 VDPWR.n543 VGND 0.100448f
C4746 VDPWR.t402 VGND 0.050988f
C4747 VDPWR.n544 VGND 0.095922f
C4748 VDPWR.n545 VGND 0.062776f
C4749 VDPWR.n546 VGND 0.037653f
C4750 VDPWR.t154 VGND 0.051359f
C4751 VDPWR.t383 VGND 0.050988f
C4752 VDPWR.n547 VGND 0.189533f
C4753 VDPWR.t576 VGND 0.050988f
C4754 VDPWR.n548 VGND 0.100448f
C4755 VDPWR.t588 VGND 0.050988f
C4756 VDPWR.n549 VGND 0.095922f
C4757 VDPWR.n550 VGND 0.271631f
C4758 VDPWR.n551 VGND 0.037653f
C4759 VDPWR.n552 VGND 0.309732f
C4760 VDPWR.n553 VGND 0.123112f
C4761 VDPWR.t153 VGND 0.669317f
C4762 VDPWR.n554 VGND 0.157342f
C4763 VDPWR.n555 VGND 0.375026f
C4764 VDPWR.n556 VGND 0.399471f
C4765 VDPWR.n557 VGND 0.042196f
C4766 VDPWR.n558 VGND 0.036863f
C4767 VDPWR.n559 VGND 0.042196f
C4768 VDPWR.n560 VGND 0.074675f
C4769 VDPWR.n561 VGND 0.046883f
C4770 VDPWR.n562 VGND 0.006668f
C4771 VDPWR.n563 VGND 0.508713f
C4772 VDPWR.n564 VGND 0.079438f
C4773 VDPWR.n565 VGND 0.079438f
C4774 VDPWR.n566 VGND 0.066601f
C4775 VDPWR.n567 VGND 0.108613f
C4776 VDPWR.n568 VGND 0.204811f
C4777 VDPWR.n569 VGND 0.151285f
C4778 VDPWR.n570 VGND 0.123112f
C4779 VDPWR.t260 VGND 0.669317f
C4780 VDPWR.n571 VGND 0.157342f
C4781 VDPWR.n572 VGND 0.375026f
C4782 VDPWR.n573 VGND 0.399471f
C4783 VDPWR.n574 VGND 0.042196f
C4784 VDPWR.n575 VGND 0.036863f
C4785 VDPWR.n576 VGND 0.042196f
C4786 VDPWR.n577 VGND 0.074675f
C4787 VDPWR.n578 VGND 0.046883f
C4788 VDPWR.n579 VGND 0.006668f
C4789 VDPWR.n580 VGND 0.508713f
C4790 VDPWR.n581 VGND 0.079438f
C4791 VDPWR.n582 VGND 0.079438f
C4792 VDPWR.n583 VGND 0.066601f
C4793 VDPWR.n584 VGND 0.108613f
C4794 VDPWR.n585 VGND 0.204811f
C4795 VDPWR.n586 VGND 0.151285f
C4796 VDPWR.n587 VGND 0.123112f
C4797 VDPWR.t246 VGND 0.669317f
C4798 VDPWR.n588 VGND 0.157342f
C4799 VDPWR.n589 VGND 0.375026f
C4800 VDPWR.n590 VGND 0.399471f
C4801 VDPWR.n591 VGND 0.042196f
C4802 VDPWR.n592 VGND 0.036863f
C4803 VDPWR.n593 VGND 0.042196f
C4804 VDPWR.n594 VGND 0.074675f
C4805 VDPWR.n595 VGND 0.046883f
C4806 VDPWR.n596 VGND 0.006668f
C4807 VDPWR.n597 VGND 0.508713f
C4808 VDPWR.n598 VGND 0.079438f
C4809 VDPWR.n599 VGND 0.079438f
C4810 VDPWR.n600 VGND 0.066601f
C4811 VDPWR.n601 VGND 0.108613f
C4812 VDPWR.n602 VGND 0.204811f
C4813 VDPWR.n603 VGND 0.151285f
C4814 VDPWR.n604 VGND 0.123112f
C4815 VDPWR.t122 VGND 0.669317f
C4816 VDPWR.n605 VGND 0.157342f
C4817 VDPWR.n606 VGND 0.375026f
C4818 VDPWR.n607 VGND 0.399471f
C4819 VDPWR.n608 VGND 0.042196f
C4820 VDPWR.n609 VGND 0.036863f
C4821 VDPWR.n610 VGND 0.042196f
C4822 VDPWR.n611 VGND 0.074675f
C4823 VDPWR.n612 VGND 0.046883f
C4824 VDPWR.n613 VGND 0.006668f
C4825 VDPWR.n614 VGND 0.508713f
C4826 VDPWR.n615 VGND 0.079438f
C4827 VDPWR.n616 VGND 0.079438f
C4828 VDPWR.n617 VGND 0.066601f
C4829 VDPWR.n618 VGND 0.108613f
C4830 VDPWR.n619 VGND 0.204811f
C4831 VDPWR.n620 VGND 0.151285f
C4832 VDPWR.n621 VGND 0.123112f
C4833 VDPWR.t186 VGND 0.669317f
C4834 VDPWR.n622 VGND 0.157342f
C4835 VDPWR.n623 VGND 0.375026f
C4836 VDPWR.n624 VGND 0.399471f
C4837 VDPWR.n625 VGND 0.042196f
C4838 VDPWR.n626 VGND 0.036863f
C4839 VDPWR.n627 VGND 0.042196f
C4840 VDPWR.n628 VGND 0.074675f
C4841 VDPWR.n629 VGND 0.046883f
C4842 VDPWR.n630 VGND 0.006668f
C4843 VDPWR.n631 VGND 0.508713f
C4844 VDPWR.n632 VGND 0.079438f
C4845 VDPWR.n633 VGND 0.079438f
C4846 VDPWR.n634 VGND 0.066601f
C4847 VDPWR.n635 VGND 0.108613f
C4848 VDPWR.n636 VGND 0.204811f
C4849 VDPWR.n637 VGND 0.151285f
C4850 VDPWR.n638 VGND 0.123112f
C4851 VDPWR.t315 VGND 0.669317f
C4852 VDPWR.n639 VGND 0.157342f
C4853 VDPWR.n640 VGND 0.375026f
C4854 VDPWR.n641 VGND 0.399471f
C4855 VDPWR.n642 VGND 0.042196f
C4856 VDPWR.n643 VGND 0.036863f
C4857 VDPWR.n644 VGND 0.042196f
C4858 VDPWR.n645 VGND 0.074675f
C4859 VDPWR.n646 VGND 0.046883f
C4860 VDPWR.n647 VGND 0.006668f
C4861 VDPWR.n648 VGND 0.508713f
C4862 VDPWR.n649 VGND 0.079438f
C4863 VDPWR.n650 VGND 0.079438f
C4864 VDPWR.n651 VGND 0.066601f
C4865 VDPWR.n652 VGND 0.108613f
C4866 VDPWR.n653 VGND 0.204811f
C4867 VDPWR.n654 VGND 0.151285f
C4868 VDPWR.n655 VGND 0.123112f
C4869 VDPWR.t214 VGND 0.669317f
C4870 VDPWR.n656 VGND 0.157342f
C4871 VDPWR.n657 VGND 0.375026f
C4872 VDPWR.n658 VGND 0.399471f
C4873 VDPWR.n659 VGND 0.042196f
C4874 VDPWR.n660 VGND 0.036863f
C4875 VDPWR.n661 VGND 0.042196f
C4876 VDPWR.n662 VGND 0.074675f
C4877 VDPWR.n663 VGND 0.046883f
C4878 VDPWR.n664 VGND 0.006668f
C4879 VDPWR.n665 VGND 0.508713f
C4880 VDPWR.n666 VGND 0.079438f
C4881 VDPWR.n667 VGND 0.079438f
C4882 VDPWR.n668 VGND 0.066601f
C4883 VDPWR.n669 VGND 0.108613f
C4884 VDPWR.n670 VGND 0.204811f
C4885 VDPWR.n671 VGND 0.151285f
C4886 VDPWR.n672 VGND 0.123112f
C4887 VDPWR.t71 VGND 0.669317f
C4888 VDPWR.n673 VGND 0.157342f
C4889 VDPWR.n674 VGND 0.375026f
C4890 VDPWR.n675 VGND 0.399471f
C4891 VDPWR.n676 VGND 0.042196f
C4892 VDPWR.n677 VGND 0.036863f
C4893 VDPWR.n678 VGND 0.042196f
C4894 VDPWR.n679 VGND 0.074675f
C4895 VDPWR.n680 VGND 0.046883f
C4896 VDPWR.n681 VGND 0.006668f
C4897 VDPWR.n682 VGND 0.508713f
C4898 VDPWR.n683 VGND 0.079438f
C4899 VDPWR.n684 VGND 0.079438f
C4900 VDPWR.n685 VGND 0.066601f
C4901 VDPWR.n686 VGND 0.108613f
C4902 VDPWR.n687 VGND 0.047195f
C4903 VDPWR.t607 VGND 0.05099f
C4904 VDPWR.n688 VGND 0.094073f
C4905 VDPWR.n689 VGND 0.041613f
C4906 VDPWR.n690 VGND 0.043998f
C4907 VDPWR.n691 VGND 0.02174f
C4908 VDPWR.n692 VGND 0.031242f
C4909 VDPWR.n693 VGND 0.052314f
C4910 VDPWR.t150 VGND 0.05099f
C4911 VDPWR.n694 VGND 0.043998f
C4912 VDPWR.t110 VGND 0.05099f
C4913 VDPWR.n695 VGND 0.094073f
C4914 VDPWR.n696 VGND 0.02174f
C4915 VDPWR.n697 VGND 0.043998f
C4916 VDPWR.n698 VGND 0.02174f
C4917 VDPWR.n699 VGND 0.031242f
C4918 VDPWR.n700 VGND 0.052314f
C4919 VDPWR.t147 VGND 0.05099f
C4920 VDPWR.n701 VGND 0.043998f
C4921 VDPWR.t405 VGND 0.05099f
C4922 VDPWR.n702 VGND 0.094073f
C4923 VDPWR.n703 VGND 0.02174f
C4924 VDPWR.n704 VGND 0.043998f
C4925 VDPWR.n705 VGND 0.02174f
C4926 VDPWR.n706 VGND 0.031242f
C4927 VDPWR.n707 VGND 0.052314f
C4928 VDPWR.t193 VGND 0.05099f
C4929 VDPWR.n708 VGND 0.043998f
C4930 VDPWR.t609 VGND 0.05099f
C4931 VDPWR.n709 VGND 0.094073f
C4932 VDPWR.n710 VGND 0.02174f
C4933 VDPWR.n711 VGND 0.043998f
C4934 VDPWR.n712 VGND 0.02174f
C4935 VDPWR.n713 VGND 0.031242f
C4936 VDPWR.n714 VGND 0.052314f
C4937 VDPWR.t404 VGND 0.05099f
C4938 VDPWR.n715 VGND 0.043998f
C4939 VDPWR.t173 VGND 0.05099f
C4940 VDPWR.n716 VGND 0.094073f
C4941 VDPWR.n717 VGND 0.02174f
C4942 VDPWR.n718 VGND 0.043998f
C4943 VDPWR.n719 VGND 0.02174f
C4944 VDPWR.n720 VGND 0.031242f
C4945 VDPWR.n721 VGND 0.052314f
C4946 VDPWR.t602 VGND 0.05099f
C4947 VDPWR.n722 VGND 0.043998f
C4948 VDPWR.t172 VGND 0.05099f
C4949 VDPWR.n723 VGND 0.094073f
C4950 VDPWR.n724 VGND 0.02174f
C4951 VDPWR.n725 VGND 0.043998f
C4952 VDPWR.n726 VGND 0.02174f
C4953 VDPWR.n727 VGND 0.031242f
C4954 VDPWR.n728 VGND 0.052314f
C4955 VDPWR.t601 VGND 0.05099f
C4956 VDPWR.n729 VGND 0.043998f
C4957 VDPWR.t192 VGND 0.05099f
C4958 VDPWR.n730 VGND 0.094073f
C4959 VDPWR.n731 VGND 0.02174f
C4960 VDPWR.n732 VGND 0.043998f
C4961 VDPWR.n733 VGND 0.02174f
C4962 VDPWR.n734 VGND 0.031242f
C4963 VDPWR.n735 VGND 0.052314f
C4964 VDPWR.t608 VGND 0.05099f
C4965 VDPWR.n736 VGND 0.043998f
C4966 VDPWR.t403 VGND 0.05099f
C4967 VDPWR.n737 VGND 0.094073f
C4968 VDPWR.n738 VGND 0.02174f
C4969 VDPWR.n739 VGND 0.043998f
C4970 VDPWR.n740 VGND 0.02174f
C4971 VDPWR.n741 VGND 0.031242f
C4972 VDPWR.n742 VGND 0.052314f
C4973 VDPWR.t111 VGND 0.05099f
C4974 VDPWR.n743 VGND 0.043998f
C4975 VDPWR.t554 VGND 0.05099f
C4976 VDPWR.n744 VGND 0.094073f
C4977 VDPWR.n745 VGND 0.02174f
C4978 VDPWR.n746 VGND 0.043998f
C4979 VDPWR.n747 VGND 0.02174f
C4980 VDPWR.n748 VGND 0.031242f
C4981 VDPWR.n749 VGND 0.052314f
C4982 VDPWR.t556 VGND 0.05099f
C4983 VDPWR.n750 VGND 0.043998f
C4984 VDPWR.t557 VGND 0.05099f
C4985 VDPWR.n751 VGND 0.094073f
C4986 VDPWR.n752 VGND 0.02174f
C4987 VDPWR.n753 VGND 0.043998f
C4988 VDPWR.n754 VGND 0.02174f
C4989 VDPWR.n755 VGND 0.031242f
C4990 VDPWR.n756 VGND 0.052314f
C4991 VDPWR.t555 VGND 0.05099f
C4992 VDPWR.n757 VGND 0.043998f
C4993 VDPWR.t25 VGND 0.05099f
C4994 VDPWR.n758 VGND 0.094073f
C4995 VDPWR.n759 VGND 0.02174f
C4996 VDPWR.n760 VGND 0.043998f
C4997 VDPWR.n761 VGND 0.02174f
C4998 VDPWR.n762 VGND 0.031242f
C4999 VDPWR.n763 VGND 0.052314f
C5000 VDPWR.t482 VGND 0.05099f
C5001 VDPWR.n764 VGND 0.043998f
C5002 VDPWR.t103 VGND 0.05099f
C5003 VDPWR.n765 VGND 0.094073f
C5004 VDPWR.n766 VGND 0.02174f
C5005 VDPWR.n767 VGND 0.043998f
C5006 VDPWR.n768 VGND 0.02174f
C5007 VDPWR.n769 VGND 0.031242f
C5008 VDPWR.n770 VGND 0.052314f
C5009 VDPWR.t594 VGND 0.05099f
C5010 VDPWR.n771 VGND 0.043998f
C5011 VDPWR.t265 VGND 0.05099f
C5012 VDPWR.n772 VGND 0.094073f
C5013 VDPWR.n773 VGND 0.02174f
C5014 VDPWR.n774 VGND 0.043998f
C5015 VDPWR.n775 VGND 0.02174f
C5016 VDPWR.n776 VGND 0.031242f
C5017 VDPWR.n777 VGND 0.052314f
C5018 VDPWR.t597 VGND 0.05099f
C5019 VDPWR.n778 VGND 0.043998f
C5020 VDPWR.t81 VGND 0.05099f
C5021 VDPWR.n779 VGND 0.094073f
C5022 VDPWR.n780 VGND 0.02174f
C5023 VDPWR.n781 VGND 0.043998f
C5024 VDPWR.n782 VGND 0.041613f
C5025 VDPWR.t24 VGND 4.806f
C5026 VDPWR.n783 VGND 0.03114f
C5027 VDPWR.n784 VGND 0.031242f
C5028 VDPWR.n785 VGND 0.027943f
C5029 VDPWR.n786 VGND 0.031242f
C5030 VDPWR.n787 VGND 0.027943f
C5031 VDPWR.n788 VGND 0.031242f
C5032 VDPWR.n789 VGND 0.027943f
C5033 VDPWR.n790 VGND 0.031242f
C5034 VDPWR.n791 VGND 0.027943f
C5035 VDPWR.n792 VGND 0.031242f
C5036 VDPWR.n793 VGND 0.027943f
C5037 VDPWR.n794 VGND 0.031242f
C5038 VDPWR.n795 VGND 0.027943f
C5039 VDPWR.n796 VGND 0.031242f
C5040 VDPWR.n797 VGND 0.027943f
C5041 VDPWR.n798 VGND 0.031242f
C5042 VDPWR.n799 VGND 0.027943f
C5043 VDPWR.n800 VGND 0.031242f
C5044 VDPWR.n801 VGND 0.027943f
C5045 VDPWR.n802 VGND 0.031242f
C5046 VDPWR.n803 VGND 0.027943f
C5047 VDPWR.n804 VGND 0.031242f
C5048 VDPWR.n805 VGND 0.027943f
C5049 VDPWR.n806 VGND 0.031242f
C5050 VDPWR.n807 VGND 0.027943f
C5051 VDPWR.n808 VGND 0.031242f
C5052 VDPWR.n809 VGND 0.027943f
C5053 VDPWR.n810 VGND 0.031242f
C5054 VDPWR.n811 VGND 0.027943f
C5055 VDPWR.n812 VGND 0.031242f
C5056 VDPWR.n813 VGND 0.027943f
C5057 VDPWR.n814 VGND 0.031242f
C5058 VDPWR.n815 VGND 0.027943f
C5059 VDPWR.n816 VGND 0.031242f
C5060 VDPWR.n817 VGND 0.027943f
C5061 VDPWR.n818 VGND 0.031242f
C5062 VDPWR.n819 VGND 0.027943f
C5063 VDPWR.n820 VGND 0.031242f
C5064 VDPWR.n821 VGND 0.027943f
C5065 VDPWR.n822 VGND 0.031242f
C5066 VDPWR.n823 VGND 0.027943f
C5067 VDPWR.n824 VGND 0.031242f
C5068 VDPWR.n825 VGND 0.027943f
C5069 VDPWR.n826 VGND 0.031242f
C5070 VDPWR.n827 VGND 0.027943f
C5071 VDPWR.n828 VGND 0.031242f
C5072 VDPWR.n829 VGND 0.027943f
C5073 VDPWR.n830 VGND 0.031242f
C5074 VDPWR.n831 VGND 0.027943f
C5075 VDPWR.n832 VGND 0.031242f
C5076 VDPWR.n833 VGND 0.027943f
C5077 VDPWR.n834 VGND 0.031242f
C5078 VDPWR.n835 VGND 0.027943f
C5079 VDPWR.n836 VGND 3.55953f
C5080 VDPWR.n837 VGND 0.031242f
C5081 VDPWR.n838 VGND 0.027943f
C5082 VDPWR.n839 VGND 2.63431f
C5083 VDPWR.n840 VGND 0.03114f
C5084 VDPWR.n841 VGND 0.047195f
C5085 VDPWR.n842 VGND 0.052314f
C5086 VDPWR.t141 VGND 0.05099f
C5087 VDPWR.n843 VGND 0.045492f
C5088 VDPWR.n844 VGND 0.094073f
C5089 VDPWR.n845 VGND 0.014168f
C5090 VDPWR.n846 VGND 0.041613f
C5091 VDPWR.n847 VGND 0.031242f
C5092 VDPWR.n848 VGND 0.02174f
C5093 VDPWR.n849 VGND 0.014168f
C5094 VDPWR.n850 VGND 0.052314f
C5095 VDPWR.n851 VGND 0.094073f
C5096 VDPWR.n852 VGND 0.014168f
C5097 VDPWR.n853 VGND 0.02174f
C5098 VDPWR.n854 VGND 0.031242f
C5099 VDPWR.n855 VGND 0.02174f
C5100 VDPWR.n856 VGND 0.014168f
C5101 VDPWR.n857 VGND 0.052314f
C5102 VDPWR.n858 VGND 0.094073f
C5103 VDPWR.n859 VGND 0.014168f
C5104 VDPWR.n860 VGND 0.02174f
C5105 VDPWR.n861 VGND 0.031242f
C5106 VDPWR.n862 VGND 0.02174f
C5107 VDPWR.n863 VGND 0.014168f
C5108 VDPWR.n864 VGND 0.052314f
C5109 VDPWR.n865 VGND 0.094073f
C5110 VDPWR.n866 VGND 0.014168f
C5111 VDPWR.n867 VGND 0.02174f
C5112 VDPWR.n868 VGND 0.031242f
C5113 VDPWR.n869 VGND 0.02174f
C5114 VDPWR.n870 VGND 0.014168f
C5115 VDPWR.n871 VGND 0.052314f
C5116 VDPWR.n872 VGND 0.094073f
C5117 VDPWR.n873 VGND 0.014168f
C5118 VDPWR.n874 VGND 0.02174f
C5119 VDPWR.n875 VGND 0.031242f
C5120 VDPWR.n876 VGND 0.02174f
C5121 VDPWR.n877 VGND 0.014168f
C5122 VDPWR.n878 VGND 0.052314f
C5123 VDPWR.n879 VGND 0.094073f
C5124 VDPWR.n880 VGND 0.014168f
C5125 VDPWR.n881 VGND 0.02174f
C5126 VDPWR.n882 VGND 0.031242f
C5127 VDPWR.n883 VGND 0.02174f
C5128 VDPWR.n884 VGND 0.014168f
C5129 VDPWR.n885 VGND 0.052314f
C5130 VDPWR.n886 VGND 0.094073f
C5131 VDPWR.n887 VGND 0.014168f
C5132 VDPWR.n888 VGND 0.02174f
C5133 VDPWR.n889 VGND 0.031242f
C5134 VDPWR.n890 VGND 0.02174f
C5135 VDPWR.n891 VGND 0.014168f
C5136 VDPWR.n892 VGND 0.052314f
C5137 VDPWR.n893 VGND 0.094073f
C5138 VDPWR.n894 VGND 0.014168f
C5139 VDPWR.n895 VGND 0.02174f
C5140 VDPWR.n896 VGND 0.031242f
C5141 VDPWR.n897 VGND 0.02174f
C5142 VDPWR.n898 VGND 0.014168f
C5143 VDPWR.n899 VGND 0.052314f
C5144 VDPWR.n900 VGND 0.094073f
C5145 VDPWR.n901 VGND 0.014168f
C5146 VDPWR.n902 VGND 0.02174f
C5147 VDPWR.n903 VGND 0.031242f
C5148 VDPWR.n904 VGND 0.02174f
C5149 VDPWR.n905 VGND 0.014168f
C5150 VDPWR.n906 VGND 0.052314f
C5151 VDPWR.n907 VGND 0.094073f
C5152 VDPWR.n908 VGND 0.014168f
C5153 VDPWR.n909 VGND 0.02174f
C5154 VDPWR.n910 VGND 0.031242f
C5155 VDPWR.n911 VGND 0.02174f
C5156 VDPWR.n912 VGND 0.014168f
C5157 VDPWR.n913 VGND 0.052314f
C5158 VDPWR.n914 VGND 0.094073f
C5159 VDPWR.n915 VGND 0.014168f
C5160 VDPWR.n916 VGND 0.02174f
C5161 VDPWR.n917 VGND 0.031242f
C5162 VDPWR.n918 VGND 0.02174f
C5163 VDPWR.n919 VGND 0.014168f
C5164 VDPWR.n920 VGND 0.052314f
C5165 VDPWR.n921 VGND 0.094073f
C5166 VDPWR.n922 VGND 0.014168f
C5167 VDPWR.n923 VGND 0.02174f
C5168 VDPWR.n924 VGND 0.031242f
C5169 VDPWR.n925 VGND 0.02174f
C5170 VDPWR.n926 VGND 0.014168f
C5171 VDPWR.n927 VGND 0.052314f
C5172 VDPWR.n928 VGND 0.094073f
C5173 VDPWR.n929 VGND 0.014168f
C5174 VDPWR.n930 VGND 0.02174f
C5175 VDPWR.n931 VGND 0.031242f
C5176 VDPWR.n932 VGND 0.02174f
C5177 VDPWR.n933 VGND 0.014168f
C5178 VDPWR.n934 VGND 0.052314f
C5179 VDPWR.n935 VGND 0.094073f
C5180 VDPWR.n936 VGND 0.014168f
C5181 VDPWR.n937 VGND 0.02174f
C5182 VDPWR.n938 VGND 0.031242f
C5183 VDPWR.n939 VGND 0.041613f
C5184 VDPWR.n940 VGND 0.014168f
C5185 VDPWR.n941 VGND 0.099317f
C5186 VDPWR.n942 VGND 0.069883f
C5187 VDPWR.t346 VGND 0.013587f
C5188 VDPWR.t600 VGND 0.013587f
C5189 VDPWR.n943 VGND 0.028793f
C5190 VDPWR.t392 VGND 0.051222f
C5191 VDPWR.n944 VGND 0.04964f
C5192 VDPWR.t389 VGND 0.051222f
C5193 VDPWR.n945 VGND 0.11792f
C5194 VDPWR.n946 VGND 0.069883f
C5195 VDPWR.t205 VGND 0.013587f
C5196 VDPWR.t587 VGND 0.013587f
C5197 VDPWR.n947 VGND 0.028793f
C5198 VDPWR.t211 VGND 0.051222f
C5199 VDPWR.n948 VGND 0.04964f
C5200 VDPWR.t263 VGND 0.051222f
C5201 VDPWR.n949 VGND 0.11792f
C5202 VDPWR.n950 VGND 0.069883f
C5203 VDPWR.t318 VGND 0.013587f
C5204 VDPWR.t325 VGND 0.013587f
C5205 VDPWR.n951 VGND 0.028793f
C5206 VDPWR.t143 VGND 0.051222f
C5207 VDPWR.n952 VGND 0.04964f
C5208 VDPWR.t105 VGND 0.051222f
C5209 VDPWR.n953 VGND 0.11792f
C5210 VDPWR.n954 VGND 0.069883f
C5211 VDPWR.t183 VGND 0.013587f
C5212 VDPWR.t156 VGND 0.013587f
C5213 VDPWR.n955 VGND 0.028793f
C5214 VDPWR.t9 VGND 0.051222f
C5215 VDPWR.n956 VGND 0.04964f
C5216 VDPWR.t382 VGND 0.051222f
C5217 VDPWR.n957 VGND 0.11792f
C5218 VDPWR.n958 VGND 0.069883f
C5219 VDPWR.t357 VGND 0.013587f
C5220 VDPWR.t238 VGND 0.013587f
C5221 VDPWR.n959 VGND 0.028793f
C5222 VDPWR.t566 VGND 0.051222f
C5223 VDPWR.n960 VGND 0.04964f
C5224 VDPWR.t522 VGND 0.051222f
C5225 VDPWR.n961 VGND 0.11792f
C5226 VDPWR.n962 VGND 0.069883f
C5227 VDPWR.t400 VGND 0.013587f
C5228 VDPWR.t249 VGND 0.013587f
C5229 VDPWR.n963 VGND 0.028793f
C5230 VDPWR.t7 VGND 0.051222f
C5231 VDPWR.n964 VGND 0.04964f
C5232 VDPWR.t280 VGND 0.051222f
C5233 VDPWR.n965 VGND 0.11792f
C5234 VDPWR.n966 VGND 0.069883f
C5235 VDPWR.t581 VGND 0.013587f
C5236 VDPWR.t168 VGND 0.013587f
C5237 VDPWR.n967 VGND 0.028793f
C5238 VDPWR.t500 VGND 0.051222f
C5239 VDPWR.n968 VGND 0.04964f
C5240 VDPWR.t494 VGND 0.051222f
C5241 VDPWR.n969 VGND 0.11792f
C5242 VDPWR.n970 VGND 0.069883f
C5243 VDPWR.t498 VGND 0.013587f
C5244 VDPWR.t578 VGND 0.013587f
C5245 VDPWR.n971 VGND 0.028793f
C5246 VDPWR.t32 VGND 0.051222f
C5247 VDPWR.n972 VGND 0.04964f
C5248 VDPWR.t218 VGND 0.051222f
C5249 VDPWR.n973 VGND 0.11792f
C5250 VDPWR.t385 VGND 0.013587f
C5251 VDPWR.t170 VGND 0.013587f
C5252 VDPWR.n974 VGND 0.028793f
C5253 VDPWR.n975 VGND 0.246742f
C5254 VDPWR.n976 VGND 0.083093f
C5255 VDPWR.n977 VGND 0.26841f
C5256 VDPWR.n978 VGND 0.101548f
C5257 VDPWR.t384 VGND 0.209173f
C5258 VDPWR.t169 VGND 0.131939f
C5259 VDPWR.t33 VGND 0.131939f
C5260 VDPWR.t217 VGND 0.173169f
C5261 VDPWR.n979 VGND 0.265912f
C5262 VDPWR.t577 VGND 0.205573f
C5263 VDPWR.t497 VGND 0.131939f
C5264 VDPWR.t128 VGND 0.131939f
C5265 VDPWR.t31 VGND 0.174669f
C5266 VDPWR.n980 VGND 0.029939f
C5267 VDPWR.n981 VGND 0.110199f
C5268 VDPWR.n982 VGND 0.108699f
C5269 VDPWR.n983 VGND 0.089537f
C5270 VDPWR.n984 VGND 0.101548f
C5271 VDPWR.n985 VGND 0.089537f
C5272 VDPWR.n986 VGND 0.008045f
C5273 VDPWR.n987 VGND 0.044727f
C5274 VDPWR.n988 VGND 0.118079f
C5275 VDPWR.n989 VGND 0.120342f
C5276 VDPWR.n990 VGND 0.058904f
C5277 VDPWR.t64 VGND 0.013587f
C5278 VDPWR.t370 VGND 0.013587f
C5279 VDPWR.n991 VGND 0.028793f
C5280 VDPWR.n992 VGND 0.12082f
C5281 VDPWR.n993 VGND 0.095544f
C5282 VDPWR.n994 VGND 0.069983f
C5283 VDPWR.n995 VGND 0.26841f
C5284 VDPWR.n996 VGND 0.101548f
C5285 VDPWR.t63 VGND 0.209173f
C5286 VDPWR.t369 VGND 0.131939f
C5287 VDPWR.t533 VGND 0.131939f
C5288 VDPWR.t493 VGND 0.173169f
C5289 VDPWR.n997 VGND 0.265912f
C5290 VDPWR.t167 VGND 0.205573f
C5291 VDPWR.t580 VGND 0.131939f
C5292 VDPWR.t245 VGND 0.131939f
C5293 VDPWR.t499 VGND 0.174669f
C5294 VDPWR.n998 VGND 0.029939f
C5295 VDPWR.n999 VGND 0.110199f
C5296 VDPWR.n1000 VGND 0.108699f
C5297 VDPWR.n1001 VGND 0.089537f
C5298 VDPWR.n1002 VGND 0.101548f
C5299 VDPWR.n1003 VGND 0.089537f
C5300 VDPWR.n1004 VGND 0.008045f
C5301 VDPWR.n1005 VGND 0.044727f
C5302 VDPWR.n1006 VGND 0.118079f
C5303 VDPWR.n1007 VGND 0.120342f
C5304 VDPWR.n1008 VGND 0.058904f
C5305 VDPWR.t398 VGND 0.013587f
C5306 VDPWR.t115 VGND 0.013587f
C5307 VDPWR.n1009 VGND 0.028793f
C5308 VDPWR.n1010 VGND 0.12082f
C5309 VDPWR.n1011 VGND 0.095544f
C5310 VDPWR.n1012 VGND 0.069983f
C5311 VDPWR.n1013 VGND 0.26841f
C5312 VDPWR.n1014 VGND 0.101548f
C5313 VDPWR.t397 VGND 0.209173f
C5314 VDPWR.t114 VGND 0.131939f
C5315 VDPWR.t266 VGND 0.131939f
C5316 VDPWR.t279 VGND 0.173169f
C5317 VDPWR.n1015 VGND 0.265912f
C5318 VDPWR.t248 VGND 0.205573f
C5319 VDPWR.t399 VGND 0.131939f
C5320 VDPWR.t510 VGND 0.131939f
C5321 VDPWR.t6 VGND 0.174669f
C5322 VDPWR.n1016 VGND 0.029939f
C5323 VDPWR.n1017 VGND 0.110199f
C5324 VDPWR.n1018 VGND 0.108699f
C5325 VDPWR.n1019 VGND 0.089537f
C5326 VDPWR.n1020 VGND 0.101548f
C5327 VDPWR.n1021 VGND 0.089537f
C5328 VDPWR.n1022 VGND 0.008045f
C5329 VDPWR.n1023 VGND 0.044727f
C5330 VDPWR.n1024 VGND 0.118079f
C5331 VDPWR.n1025 VGND 0.120342f
C5332 VDPWR.n1026 VGND 0.058904f
C5333 VDPWR.t146 VGND 0.013587f
C5334 VDPWR.t236 VGND 0.013587f
C5335 VDPWR.n1027 VGND 0.028793f
C5336 VDPWR.n1028 VGND 0.12082f
C5337 VDPWR.n1029 VGND 0.095544f
C5338 VDPWR.n1030 VGND 0.069983f
C5339 VDPWR.n1031 VGND 0.26841f
C5340 VDPWR.n1032 VGND 0.101548f
C5341 VDPWR.t145 VGND 0.209173f
C5342 VDPWR.t235 VGND 0.131939f
C5343 VDPWR.t264 VGND 0.131939f
C5344 VDPWR.t521 VGND 0.173169f
C5345 VDPWR.n1033 VGND 0.265912f
C5346 VDPWR.t237 VGND 0.205573f
C5347 VDPWR.t356 VGND 0.131939f
C5348 VDPWR.t28 VGND 0.131939f
C5349 VDPWR.t565 VGND 0.174669f
C5350 VDPWR.n1034 VGND 0.029939f
C5351 VDPWR.n1035 VGND 0.110199f
C5352 VDPWR.n1036 VGND 0.108699f
C5353 VDPWR.n1037 VGND 0.089537f
C5354 VDPWR.n1038 VGND 0.101548f
C5355 VDPWR.n1039 VGND 0.089537f
C5356 VDPWR.n1040 VGND 0.008045f
C5357 VDPWR.n1041 VGND 0.044727f
C5358 VDPWR.n1042 VGND 0.118079f
C5359 VDPWR.n1043 VGND 0.120342f
C5360 VDPWR.n1044 VGND 0.058904f
C5361 VDPWR.t185 VGND 0.013587f
C5362 VDPWR.t362 VGND 0.013587f
C5363 VDPWR.n1045 VGND 0.028793f
C5364 VDPWR.n1046 VGND 0.12082f
C5365 VDPWR.n1047 VGND 0.095544f
C5366 VDPWR.n1048 VGND 0.069983f
C5367 VDPWR.n1049 VGND 0.26841f
C5368 VDPWR.n1050 VGND 0.101548f
C5369 VDPWR.t184 VGND 0.209173f
C5370 VDPWR.t361 VGND 0.131939f
C5371 VDPWR.t84 VGND 0.131939f
C5372 VDPWR.t381 VGND 0.173169f
C5373 VDPWR.n1051 VGND 0.265912f
C5374 VDPWR.t155 VGND 0.205573f
C5375 VDPWR.t182 VGND 0.131939f
C5376 VDPWR.t596 VGND 0.131939f
C5377 VDPWR.t8 VGND 0.174669f
C5378 VDPWR.n1052 VGND 0.029939f
C5379 VDPWR.n1053 VGND 0.110199f
C5380 VDPWR.n1054 VGND 0.108699f
C5381 VDPWR.n1055 VGND 0.089537f
C5382 VDPWR.n1056 VGND 0.101548f
C5383 VDPWR.n1057 VGND 0.089537f
C5384 VDPWR.n1058 VGND 0.008045f
C5385 VDPWR.n1059 VGND 0.044727f
C5386 VDPWR.n1060 VGND 0.118079f
C5387 VDPWR.n1061 VGND 0.120342f
C5388 VDPWR.n1062 VGND 0.058904f
C5389 VDPWR.t320 VGND 0.013587f
C5390 VDPWR.t323 VGND 0.013587f
C5391 VDPWR.n1063 VGND 0.028793f
C5392 VDPWR.n1064 VGND 0.12082f
C5393 VDPWR.n1065 VGND 0.095544f
C5394 VDPWR.n1066 VGND 0.069983f
C5395 VDPWR.n1067 VGND 0.26841f
C5396 VDPWR.n1068 VGND 0.101548f
C5397 VDPWR.t319 VGND 0.209173f
C5398 VDPWR.t322 VGND 0.131939f
C5399 VDPWR.t125 VGND 0.131939f
C5400 VDPWR.t104 VGND 0.173169f
C5401 VDPWR.n1069 VGND 0.265912f
C5402 VDPWR.t324 VGND 0.205573f
C5403 VDPWR.t317 VGND 0.131939f
C5404 VDPWR.t595 VGND 0.131939f
C5405 VDPWR.t142 VGND 0.174669f
C5406 VDPWR.n1070 VGND 0.029939f
C5407 VDPWR.n1071 VGND 0.110199f
C5408 VDPWR.n1072 VGND 0.108699f
C5409 VDPWR.n1073 VGND 0.089537f
C5410 VDPWR.n1074 VGND 0.101548f
C5411 VDPWR.n1075 VGND 0.089537f
C5412 VDPWR.n1076 VGND 0.008045f
C5413 VDPWR.n1077 VGND 0.044727f
C5414 VDPWR.n1078 VGND 0.118079f
C5415 VDPWR.n1079 VGND 0.120342f
C5416 VDPWR.n1080 VGND 0.058904f
C5417 VDPWR.t203 VGND 0.013587f
C5418 VDPWR.t425 VGND 0.013587f
C5419 VDPWR.n1081 VGND 0.028793f
C5420 VDPWR.n1082 VGND 0.12082f
C5421 VDPWR.n1083 VGND 0.095544f
C5422 VDPWR.n1084 VGND 0.069983f
C5423 VDPWR.n1085 VGND 0.26841f
C5424 VDPWR.n1086 VGND 0.101548f
C5425 VDPWR.t202 VGND 0.209173f
C5426 VDPWR.t424 VGND 0.131939f
C5427 VDPWR.t101 VGND 0.131939f
C5428 VDPWR.t262 VGND 0.173169f
C5429 VDPWR.n1087 VGND 0.265912f
C5430 VDPWR.t586 VGND 0.205573f
C5431 VDPWR.t204 VGND 0.131939f
C5432 VDPWR.t34 VGND 0.131939f
C5433 VDPWR.t210 VGND 0.174669f
C5434 VDPWR.n1088 VGND 0.029939f
C5435 VDPWR.n1089 VGND 0.110199f
C5436 VDPWR.n1090 VGND 0.108699f
C5437 VDPWR.n1091 VGND 0.089537f
C5438 VDPWR.n1092 VGND 0.101548f
C5439 VDPWR.n1093 VGND 0.089537f
C5440 VDPWR.n1094 VGND 0.008045f
C5441 VDPWR.n1095 VGND 0.044727f
C5442 VDPWR.n1096 VGND 0.118079f
C5443 VDPWR.n1097 VGND 0.120342f
C5444 VDPWR.n1098 VGND 0.058904f
C5445 VDPWR.t274 VGND 0.013587f
C5446 VDPWR.t70 VGND 0.013587f
C5447 VDPWR.n1099 VGND 0.028793f
C5448 VDPWR.n1100 VGND 0.12082f
C5449 VDPWR.n1101 VGND 0.095544f
C5450 VDPWR.n1102 VGND 0.069983f
C5451 VDPWR.n1103 VGND 0.26841f
C5452 VDPWR.n1104 VGND 0.101548f
C5453 VDPWR.t273 VGND 0.209173f
C5454 VDPWR.t69 VGND 0.131939f
C5455 VDPWR.t468 VGND 0.131939f
C5456 VDPWR.t388 VGND 0.173169f
C5457 VDPWR.n1105 VGND 0.265912f
C5458 VDPWR.t599 VGND 0.205573f
C5459 VDPWR.t345 VGND 0.131939f
C5460 VDPWR.t2 VGND 0.131939f
C5461 VDPWR.t391 VGND 0.174669f
C5462 VDPWR.n1106 VGND 0.029939f
C5463 VDPWR.n1107 VGND 0.110199f
C5464 VDPWR.n1108 VGND 0.108699f
C5465 VDPWR.n1109 VGND 0.089537f
C5466 VDPWR.n1110 VGND 0.101548f
C5467 VDPWR.n1111 VGND 0.089537f
C5468 VDPWR.n1112 VGND 0.008045f
C5469 VDPWR.n1113 VGND 0.044727f
C5470 VDPWR.n1114 VGND 0.118079f
C5471 VDPWR.n1115 VGND 0.120342f
C5472 VDPWR.n1116 VGND 0.058904f
C5473 VDPWR.n1117 VGND 0.549702f
C5474 VDPWR.n1118 VGND 0.32216f
C5475 VDPWR.n1119 VGND 0.078774f
C5476 VDPWR.t66 VGND 0.013587f
C5477 VDPWR.t225 VGND 0.013587f
C5478 VDPWR.n1120 VGND 0.029044f
C5479 VDPWR.t342 VGND 0.013587f
C5480 VDPWR.t268 VGND 0.013587f
C5481 VDPWR.n1121 VGND 0.029044f
C5482 VDPWR.t11 VGND 0.013587f
C5483 VDPWR.t5 VGND 0.013587f
C5484 VDPWR.n1122 VGND 0.029044f
C5485 VDPWR.n1123 VGND 0.117495f
C5486 VDPWR.n1124 VGND 0.078774f
C5487 VDPWR.t614 VGND 0.013587f
C5488 VDPWR.t44 VGND 0.013587f
C5489 VDPWR.n1125 VGND 0.029044f
C5490 VDPWR.t46 VGND 0.013587f
C5491 VDPWR.t529 VGND 0.013587f
C5492 VDPWR.n1126 VGND 0.029044f
C5493 VDPWR.t429 VGND 0.013587f
C5494 VDPWR.t107 VGND 0.013587f
C5495 VDPWR.n1127 VGND 0.029044f
C5496 VDPWR.n1128 VGND 0.117495f
C5497 VDPWR.n1129 VGND 0.078774f
C5498 VDPWR.t431 VGND 0.013587f
C5499 VDPWR.t409 VGND 0.013587f
C5500 VDPWR.n1130 VGND 0.029044f
C5501 VDPWR.t407 VGND 0.013587f
C5502 VDPWR.t411 VGND 0.013587f
C5503 VDPWR.n1131 VGND 0.029044f
C5504 VDPWR.t60 VGND 0.013587f
C5505 VDPWR.t58 VGND 0.013587f
C5506 VDPWR.n1132 VGND 0.029044f
C5507 VDPWR.n1133 VGND 0.117495f
C5508 VDPWR.n1134 VGND 0.078774f
C5509 VDPWR.t296 VGND 0.013587f
C5510 VDPWR.t394 VGND 0.013587f
C5511 VDPWR.n1135 VGND 0.029044f
C5512 VDPWR.t604 VGND 0.013587f
C5513 VDPWR.t396 VGND 0.013587f
C5514 VDPWR.n1136 VGND 0.029044f
C5515 VDPWR.t290 VGND 0.013587f
C5516 VDPWR.t292 VGND 0.013587f
C5517 VDPWR.n1137 VGND 0.029044f
C5518 VDPWR.n1138 VGND 0.117495f
C5519 VDPWR.n1139 VGND 0.078774f
C5520 VDPWR.t298 VGND 0.013587f
C5521 VDPWR.t484 VGND 0.013587f
C5522 VDPWR.n1140 VGND 0.029044f
C5523 VDPWR.t477 VGND 0.013587f
C5524 VDPWR.t475 VGND 0.013587f
C5525 VDPWR.n1141 VGND 0.029044f
C5526 VDPWR.t191 VGND 0.013587f
C5527 VDPWR.t189 VGND 0.013587f
C5528 VDPWR.n1142 VGND 0.029044f
C5529 VDPWR.n1143 VGND 0.117495f
C5530 VDPWR.n1144 VGND 0.078774f
C5531 VDPWR.t80 VGND 0.013587f
C5532 VDPWR.t68 VGND 0.013587f
C5533 VDPWR.n1145 VGND 0.029044f
C5534 VDPWR.t48 VGND 0.013587f
C5535 VDPWR.t496 VGND 0.013587f
C5536 VDPWR.n1146 VGND 0.029044f
C5537 VDPWR.t232 VGND 0.013587f
C5538 VDPWR.t86 VGND 0.013587f
C5539 VDPWR.n1147 VGND 0.029044f
C5540 VDPWR.n1148 VGND 0.117495f
C5541 VDPWR.n1149 VGND 0.078774f
C5542 VDPWR.t310 VGND 0.013587f
C5543 VDPWR.t257 VGND 0.013587f
C5544 VDPWR.n1150 VGND 0.029044f
C5545 VDPWR.t255 VGND 0.013587f
C5546 VDPWR.t312 VGND 0.013587f
C5547 VDPWR.n1151 VGND 0.029044f
C5548 VDPWR.t377 VGND 0.013587f
C5549 VDPWR.t240 VGND 0.013587f
C5550 VDPWR.n1152 VGND 0.029044f
C5551 VDPWR.n1153 VGND 0.117495f
C5552 VDPWR.n1154 VGND 0.078774f
C5553 VDPWR.t524 VGND 0.013587f
C5554 VDPWR.t364 VGND 0.013587f
C5555 VDPWR.n1155 VGND 0.029044f
C5556 VDPWR.t571 VGND 0.013587f
C5557 VDPWR.t569 VGND 0.013587f
C5558 VDPWR.n1156 VGND 0.029044f
C5559 VDPWR.t550 VGND 0.013587f
C5560 VDPWR.t278 VGND 0.013587f
C5561 VDPWR.n1157 VGND 0.029044f
C5562 VDPWR.n1158 VGND 0.117495f
C5563 VDPWR.n1159 VGND 0.079477f
C5564 VDPWR.t349 VGND 0.013587f
C5565 VDPWR.t177 VGND 0.013587f
C5566 VDPWR.n1160 VGND 0.029044f
C5567 VDPWR.t175 VGND 0.013587f
C5568 VDPWR.t36 VGND 0.013587f
C5569 VDPWR.n1161 VGND 0.029044f
C5570 VDPWR.t133 VGND 0.013587f
C5571 VDPWR.t228 VGND 0.013587f
C5572 VDPWR.n1162 VGND 0.029044f
C5573 VDPWR.n1163 VGND 0.117495f
C5574 VDPWR.n1164 VGND 0.095797f
C5575 VDPWR.n1165 VGND 0.091888f
C5576 VDPWR.n1166 VGND 0.053262f
C5577 VDPWR.t471 VGND 0.013587f
C5578 VDPWR.t536 VGND 0.013587f
C5579 VDPWR.n1167 VGND 0.029044f
C5580 VDPWR.n1168 VGND 0.168829f
C5581 VDPWR.n1169 VGND 0.086228f
C5582 VDPWR.n1170 VGND 0.23265f
C5583 VDPWR.t470 VGND 0.207902f
C5584 VDPWR.t535 VGND 0.140185f
C5585 VDPWR.t132 VGND 0.140185f
C5586 VDPWR.t227 VGND 0.186382f
C5587 VDPWR.n1171 VGND 0.069681f
C5588 VDPWR.n1172 VGND 0.119476f
C5589 VDPWR.n1173 VGND 0.158504f
C5590 VDPWR.t176 VGND 0.185586f
C5591 VDPWR.t348 VGND 0.140185f
C5592 VDPWR.t35 VGND 0.140185f
C5593 VDPWR.t174 VGND 0.183196f
C5594 VDPWR.n1174 VGND 0.11629f
C5595 VDPWR.n1175 VGND 0.079014f
C5596 VDPWR.n1176 VGND 0.079014f
C5597 VDPWR.n1177 VGND 0.028487f
C5598 VDPWR.n1178 VGND 0.116895f
C5599 VDPWR.n1179 VGND 0.11712f
C5600 VDPWR.n1180 VGND 0.138034f
C5601 VDPWR.t548 VGND 0.013587f
C5602 VDPWR.t552 VGND 0.013587f
C5603 VDPWR.n1181 VGND 0.029044f
C5604 VDPWR.n1182 VGND 0.11712f
C5605 VDPWR.n1183 VGND 0.138034f
C5606 VDPWR.n1184 VGND 0.078464f
C5607 VDPWR.n1185 VGND 0.171382f
C5608 VDPWR.n1186 VGND 0.231448f
C5609 VDPWR.t547 VGND 0.207902f
C5610 VDPWR.t551 VGND 0.140185f
C5611 VDPWR.t549 VGND 0.140185f
C5612 VDPWR.t277 VGND 0.186382f
C5613 VDPWR.n1187 VGND 0.052559f
C5614 VDPWR.n1188 VGND 0.158504f
C5615 VDPWR.t363 VGND 0.185586f
C5616 VDPWR.t523 VGND 0.140185f
C5617 VDPWR.t568 VGND 0.140185f
C5618 VDPWR.t570 VGND 0.183196f
C5619 VDPWR.n1189 VGND 0.11629f
C5620 VDPWR.n1190 VGND 0.185107f
C5621 VDPWR.n1191 VGND 0.007123f
C5622 VDPWR.n1192 VGND 0.175066f
C5623 VDPWR.n1193 VGND 0.028487f
C5624 VDPWR.n1194 VGND 0.116895f
C5625 VDPWR.n1195 VGND 0.11712f
C5626 VDPWR.n1196 VGND 0.138034f
C5627 VDPWR.t195 VGND 0.013587f
C5628 VDPWR.t517 VGND 0.013587f
C5629 VDPWR.n1197 VGND 0.029044f
C5630 VDPWR.n1198 VGND 0.11712f
C5631 VDPWR.n1199 VGND 0.138034f
C5632 VDPWR.n1200 VGND 0.078464f
C5633 VDPWR.n1201 VGND 0.171382f
C5634 VDPWR.n1202 VGND 0.231448f
C5635 VDPWR.t194 VGND 0.207902f
C5636 VDPWR.t516 VGND 0.140185f
C5637 VDPWR.t376 VGND 0.140185f
C5638 VDPWR.t239 VGND 0.186382f
C5639 VDPWR.n1203 VGND 0.052559f
C5640 VDPWR.n1204 VGND 0.158504f
C5641 VDPWR.t256 VGND 0.185586f
C5642 VDPWR.t309 VGND 0.140185f
C5643 VDPWR.t311 VGND 0.140185f
C5644 VDPWR.t254 VGND 0.183196f
C5645 VDPWR.n1205 VGND 0.11629f
C5646 VDPWR.n1206 VGND 0.185107f
C5647 VDPWR.n1207 VGND 0.007123f
C5648 VDPWR.n1208 VGND 0.175066f
C5649 VDPWR.n1209 VGND 0.028487f
C5650 VDPWR.n1210 VGND 0.116895f
C5651 VDPWR.n1211 VGND 0.11712f
C5652 VDPWR.n1212 VGND 0.138034f
C5653 VDPWR.t62 VGND 0.013587f
C5654 VDPWR.t538 VGND 0.013587f
C5655 VDPWR.n1213 VGND 0.029044f
C5656 VDPWR.n1214 VGND 0.11712f
C5657 VDPWR.n1215 VGND 0.138034f
C5658 VDPWR.n1216 VGND 0.078464f
C5659 VDPWR.n1217 VGND 0.171382f
C5660 VDPWR.n1218 VGND 0.231448f
C5661 VDPWR.t61 VGND 0.207902f
C5662 VDPWR.t537 VGND 0.140185f
C5663 VDPWR.t231 VGND 0.140185f
C5664 VDPWR.t85 VGND 0.186382f
C5665 VDPWR.n1219 VGND 0.052559f
C5666 VDPWR.n1220 VGND 0.158504f
C5667 VDPWR.t67 VGND 0.185586f
C5668 VDPWR.t79 VGND 0.140185f
C5669 VDPWR.t495 VGND 0.140185f
C5670 VDPWR.t47 VGND 0.183196f
C5671 VDPWR.n1221 VGND 0.11629f
C5672 VDPWR.n1222 VGND 0.185107f
C5673 VDPWR.n1223 VGND 0.007123f
C5674 VDPWR.n1224 VGND 0.175066f
C5675 VDPWR.n1225 VGND 0.028487f
C5676 VDPWR.n1226 VGND 0.116895f
C5677 VDPWR.n1227 VGND 0.11712f
C5678 VDPWR.n1228 VGND 0.138034f
C5679 VDPWR.t282 VGND 0.013587f
C5680 VDPWR.t42 VGND 0.013587f
C5681 VDPWR.n1229 VGND 0.029044f
C5682 VDPWR.n1230 VGND 0.11712f
C5683 VDPWR.n1231 VGND 0.138034f
C5684 VDPWR.n1232 VGND 0.078464f
C5685 VDPWR.n1233 VGND 0.171382f
C5686 VDPWR.n1234 VGND 0.231448f
C5687 VDPWR.t281 VGND 0.207902f
C5688 VDPWR.t41 VGND 0.140185f
C5689 VDPWR.t190 VGND 0.140185f
C5690 VDPWR.t188 VGND 0.186382f
C5691 VDPWR.n1235 VGND 0.052559f
C5692 VDPWR.n1236 VGND 0.158504f
C5693 VDPWR.t483 VGND 0.185586f
C5694 VDPWR.t297 VGND 0.140185f
C5695 VDPWR.t474 VGND 0.140185f
C5696 VDPWR.t476 VGND 0.183196f
C5697 VDPWR.n1237 VGND 0.11629f
C5698 VDPWR.n1238 VGND 0.185107f
C5699 VDPWR.n1239 VGND 0.007123f
C5700 VDPWR.n1240 VGND 0.175066f
C5701 VDPWR.n1241 VGND 0.028487f
C5702 VDPWR.n1242 VGND 0.116895f
C5703 VDPWR.n1243 VGND 0.11712f
C5704 VDPWR.n1244 VGND 0.138034f
C5705 VDPWR.t294 VGND 0.013587f
C5706 VDPWR.t288 VGND 0.013587f
C5707 VDPWR.n1245 VGND 0.029044f
C5708 VDPWR.n1246 VGND 0.11712f
C5709 VDPWR.n1247 VGND 0.138034f
C5710 VDPWR.n1248 VGND 0.078464f
C5711 VDPWR.n1249 VGND 0.171382f
C5712 VDPWR.n1250 VGND 0.231448f
C5713 VDPWR.t293 VGND 0.207902f
C5714 VDPWR.t287 VGND 0.140185f
C5715 VDPWR.t289 VGND 0.140185f
C5716 VDPWR.t291 VGND 0.186382f
C5717 VDPWR.n1251 VGND 0.052559f
C5718 VDPWR.n1252 VGND 0.158504f
C5719 VDPWR.t393 VGND 0.185586f
C5720 VDPWR.t295 VGND 0.140185f
C5721 VDPWR.t395 VGND 0.140185f
C5722 VDPWR.t603 VGND 0.183196f
C5723 VDPWR.n1253 VGND 0.11629f
C5724 VDPWR.n1254 VGND 0.185107f
C5725 VDPWR.n1255 VGND 0.007123f
C5726 VDPWR.n1256 VGND 0.175066f
C5727 VDPWR.n1257 VGND 0.028487f
C5728 VDPWR.n1258 VGND 0.116895f
C5729 VDPWR.n1259 VGND 0.11712f
C5730 VDPWR.n1260 VGND 0.138034f
C5731 VDPWR.t527 VGND 0.013587f
C5732 VDPWR.t119 VGND 0.013587f
C5733 VDPWR.n1261 VGND 0.029044f
C5734 VDPWR.n1262 VGND 0.11712f
C5735 VDPWR.n1263 VGND 0.138034f
C5736 VDPWR.n1264 VGND 0.078464f
C5737 VDPWR.n1265 VGND 0.171382f
C5738 VDPWR.n1266 VGND 0.231448f
C5739 VDPWR.t526 VGND 0.207902f
C5740 VDPWR.t118 VGND 0.140185f
C5741 VDPWR.t59 VGND 0.140185f
C5742 VDPWR.t57 VGND 0.186382f
C5743 VDPWR.n1267 VGND 0.052559f
C5744 VDPWR.n1268 VGND 0.158504f
C5745 VDPWR.t408 VGND 0.185586f
C5746 VDPWR.t430 VGND 0.140185f
C5747 VDPWR.t410 VGND 0.140185f
C5748 VDPWR.t406 VGND 0.183196f
C5749 VDPWR.n1269 VGND 0.11629f
C5750 VDPWR.n1270 VGND 0.185107f
C5751 VDPWR.n1271 VGND 0.007123f
C5752 VDPWR.n1272 VGND 0.175066f
C5753 VDPWR.n1273 VGND 0.028487f
C5754 VDPWR.n1274 VGND 0.116895f
C5755 VDPWR.n1275 VGND 0.11712f
C5756 VDPWR.n1276 VGND 0.138034f
C5757 VDPWR.t109 VGND 0.013587f
C5758 VDPWR.t38 VGND 0.013587f
C5759 VDPWR.n1277 VGND 0.029044f
C5760 VDPWR.n1278 VGND 0.11712f
C5761 VDPWR.n1279 VGND 0.138034f
C5762 VDPWR.n1280 VGND 0.078464f
C5763 VDPWR.n1281 VGND 0.171382f
C5764 VDPWR.n1282 VGND 0.231448f
C5765 VDPWR.t108 VGND 0.207902f
C5766 VDPWR.t37 VGND 0.140185f
C5767 VDPWR.t428 VGND 0.140185f
C5768 VDPWR.t106 VGND 0.186382f
C5769 VDPWR.n1283 VGND 0.052559f
C5770 VDPWR.n1284 VGND 0.158504f
C5771 VDPWR.t43 VGND 0.185586f
C5772 VDPWR.t613 VGND 0.140185f
C5773 VDPWR.t528 VGND 0.140185f
C5774 VDPWR.t45 VGND 0.183196f
C5775 VDPWR.n1285 VGND 0.11629f
C5776 VDPWR.n1286 VGND 0.185107f
C5777 VDPWR.n1287 VGND 0.007123f
C5778 VDPWR.n1288 VGND 0.175066f
C5779 VDPWR.n1289 VGND 0.028487f
C5780 VDPWR.n1290 VGND 0.116895f
C5781 VDPWR.n1291 VGND 0.11712f
C5782 VDPWR.n1292 VGND 0.138034f
C5783 VDPWR.t13 VGND 0.013587f
C5784 VDPWR.t564 VGND 0.013587f
C5785 VDPWR.n1293 VGND 0.029044f
C5786 VDPWR.n1294 VGND 0.11712f
C5787 VDPWR.n1295 VGND 0.138034f
C5788 VDPWR.n1296 VGND 0.078464f
C5789 VDPWR.n1297 VGND 0.171382f
C5790 VDPWR.n1298 VGND 0.231448f
C5791 VDPWR.t12 VGND 0.207902f
C5792 VDPWR.t563 VGND 0.140185f
C5793 VDPWR.t10 VGND 0.140185f
C5794 VDPWR.t4 VGND 0.186382f
C5795 VDPWR.n1299 VGND 0.052559f
C5796 VDPWR.n1300 VGND 0.158504f
C5797 VDPWR.t224 VGND 0.185586f
C5798 VDPWR.t65 VGND 0.140185f
C5799 VDPWR.t267 VGND 0.140185f
C5800 VDPWR.t341 VGND 0.183196f
C5801 VDPWR.n1301 VGND 0.11629f
C5802 VDPWR.n1302 VGND 0.185107f
C5803 VDPWR.n1303 VGND 0.007123f
C5804 VDPWR.n1304 VGND 0.175066f
C5805 VDPWR.n1305 VGND 0.028487f
C5806 VDPWR.n1306 VGND 0.116895f
C5807 VDPWR.n1307 VGND 0.11712f
C5808 VDPWR.n1308 VGND 0.096953f
C5809 VDPWR.n1309 VGND 0.230818f
C5810 VDPWR.n1310 VGND 6.61925f
C5811 VDPWR.n1311 VGND 0.078774f
C5812 VDPWR.t201 VGND 0.013587f
C5813 VDPWR.t230 VGND 0.013587f
C5814 VDPWR.n1312 VGND 0.029044f
C5815 VDPWR.t506 VGND 0.013587f
C5816 VDPWR.t50 VGND 0.013587f
C5817 VDPWR.n1313 VGND 0.029044f
C5818 VDPWR.t421 VGND 0.013587f
C5819 VDPWR.t300 VGND 0.013587f
C5820 VDPWR.n1314 VGND 0.029044f
C5821 VDPWR.n1315 VGND 0.117495f
C5822 VDPWR.n1316 VGND 0.078464f
C5823 VDPWR.n1317 VGND 0.171382f
C5824 VDPWR.t414 VGND 0.185586f
C5825 VDPWR.n1318 VGND 0.171693f
C5826 VDPWR.t54 VGND 0.013587f
C5827 VDPWR.t423 VGND 0.013587f
C5828 VDPWR.n1319 VGND 0.029044f
C5829 VDPWR.n1320 VGND 0.11712f
C5830 VDPWR.n1321 VGND 0.062919f
C5831 VDPWR.n1322 VGND 0.062919f
C5832 VDPWR.n1323 VGND 0.078464f
C5833 VDPWR.n1324 VGND 0.007123f
C5834 VDPWR.t74 VGND 0.013587f
C5835 VDPWR.t127 VGND 0.013587f
C5836 VDPWR.n1325 VGND 0.029044f
C5837 VDPWR.t88 VGND 0.013587f
C5838 VDPWR.t366 VGND 0.013587f
C5839 VDPWR.n1326 VGND 0.029044f
C5840 VDPWR.n1327 VGND 0.078464f
C5841 VDPWR.t314 VGND 0.013587f
C5842 VDPWR.t213 VGND 0.013587f
C5843 VDPWR.n1328 VGND 0.029044f
C5844 VDPWR.t40 VGND 0.013587f
C5845 VDPWR.t96 VGND 0.013587f
C5846 VDPWR.n1329 VGND 0.029044f
C5847 VDPWR.t344 VGND 0.013587f
C5848 VDPWR.t276 VGND 0.013587f
C5849 VDPWR.n1330 VGND 0.029044f
C5850 VDPWR.n1331 VGND 0.117495f
C5851 VDPWR.n1332 VGND 0.078464f
C5852 VDPWR.n1333 VGND 0.171693f
C5853 VDPWR.t379 VGND 0.185586f
C5854 VDPWR.n1334 VGND 0.171693f
C5855 VDPWR.t585 VGND 0.013587f
C5856 VDPWR.t272 VGND 0.013587f
C5857 VDPWR.n1335 VGND 0.029044f
C5858 VDPWR.n1336 VGND 0.11712f
C5859 VDPWR.n1337 VGND 0.062919f
C5860 VDPWR.n1338 VGND 0.062919f
C5861 VDPWR.n1339 VGND 0.078464f
C5862 VDPWR.n1340 VGND 0.007123f
C5863 VDPWR.t76 VGND 0.013587f
C5864 VDPWR.t519 VGND 0.013587f
C5865 VDPWR.n1341 VGND 0.029044f
C5866 VDPWR.t375 VGND 0.013587f
C5867 VDPWR.t531 VGND 0.013587f
C5868 VDPWR.n1342 VGND 0.029044f
C5869 VDPWR.n1343 VGND 0.078464f
C5870 VDPWR.t152 VGND 0.013587f
C5871 VDPWR.t121 VGND 0.013587f
C5872 VDPWR.n1344 VGND 0.029044f
C5873 VDPWR.t542 VGND 0.013587f
C5874 VDPWR.t158 VGND 0.013587f
C5875 VDPWR.n1345 VGND 0.029044f
C5876 VDPWR.t481 VGND 0.013587f
C5877 VDPWR.t353 VGND 0.013587f
C5878 VDPWR.n1346 VGND 0.029044f
C5879 VDPWR.n1347 VGND 0.117495f
C5880 VDPWR.n1348 VGND 0.078464f
C5881 VDPWR.n1349 VGND 0.171693f
C5882 VDPWR.t539 VGND 0.185586f
C5883 VDPWR.n1350 VGND 0.171693f
C5884 VDPWR.t351 VGND 0.013587f
C5885 VDPWR.t487 VGND 0.013587f
C5886 VDPWR.n1351 VGND 0.029044f
C5887 VDPWR.n1352 VGND 0.11712f
C5888 VDPWR.n1353 VGND 0.062919f
C5889 VDPWR.n1354 VGND 0.062919f
C5890 VDPWR.n1355 VGND 0.078464f
C5891 VDPWR.n1356 VGND 0.007123f
C5892 VDPWR.t253 VGND 0.013587f
C5893 VDPWR.t544 VGND 0.013587f
C5894 VDPWR.n1357 VGND 0.029044f
C5895 VDPWR.t546 VGND 0.013587f
C5896 VDPWR.t270 VGND 0.013587f
C5897 VDPWR.n1358 VGND 0.029044f
C5898 VDPWR.n1359 VGND 0.079477f
C5899 VDPWR.t359 VGND 0.013587f
C5900 VDPWR.t181 VGND 0.013587f
C5901 VDPWR.n1360 VGND 0.029044f
C5902 VDPWR.t575 VGND 0.013587f
C5903 VDPWR.t52 VGND 0.013587f
C5904 VDPWR.n1361 VGND 0.029044f
C5905 VDPWR.t19 VGND 0.013587f
C5906 VDPWR.t17 VGND 0.013587f
C5907 VDPWR.n1362 VGND 0.029044f
C5908 VDPWR.n1363 VGND 0.11577f
C5909 VDPWR.n1364 VGND 0.095797f
C5910 VDPWR.n1365 VGND 0.091888f
C5911 VDPWR.n1366 VGND 0.053262f
C5912 VDPWR.t15 VGND 0.013587f
C5913 VDPWR.t94 VGND 0.013587f
C5914 VDPWR.n1367 VGND 0.029201f
C5915 VDPWR.n1368 VGND 0.118612f
C5916 VDPWR.n1369 VGND 0.061604f
C5917 VDPWR.n1370 VGND 0.081955f
C5918 VDPWR.n1371 VGND 0.23265f
C5919 VDPWR.t14 VGND 0.207902f
C5920 VDPWR.t93 VGND 0.140185f
C5921 VDPWR.t18 VGND 0.140185f
C5922 VDPWR.t16 VGND 0.186382f
C5923 VDPWR.n1372 VGND 0.069681f
C5924 VDPWR.n1373 VGND 0.119476f
C5925 VDPWR.t116 VGND 0.140185f
C5926 VDPWR.t55 VGND 0.140185f
C5927 VDPWR.t233 VGND 0.183196f
C5928 VDPWR.n1374 VGND 0.11629f
C5929 VDPWR.n1375 VGND 0.185107f
C5930 VDPWR.t543 VGND 0.186382f
C5931 VDPWR.t252 VGND 0.140185f
C5932 VDPWR.t269 VGND 0.140185f
C5933 VDPWR.t545 VGND 0.185586f
C5934 VDPWR.n1376 VGND 0.052249f
C5935 VDPWR.n1377 VGND 0.207888f
C5936 VDPWR.n1378 VGND 0.158504f
C5937 VDPWR.t180 VGND 0.185586f
C5938 VDPWR.t358 VGND 0.140185f
C5939 VDPWR.t51 VGND 0.140185f
C5940 VDPWR.t574 VGND 0.183196f
C5941 VDPWR.n1379 VGND 0.11629f
C5942 VDPWR.n1380 VGND 0.079014f
C5943 VDPWR.n1381 VGND 0.079014f
C5944 VDPWR.n1382 VGND 0.028487f
C5945 VDPWR.n1383 VGND 0.116895f
C5946 VDPWR.n1384 VGND 0.11712f
C5947 VDPWR.n1385 VGND 0.062919f
C5948 VDPWR.n1386 VGND 0.062919f
C5949 VDPWR.n1387 VGND 0.11712f
C5950 VDPWR.n1388 VGND 0.117495f
C5951 VDPWR.t234 VGND 0.013587f
C5952 VDPWR.t56 VGND 0.013587f
C5953 VDPWR.n1389 VGND 0.029044f
C5954 VDPWR.t117 VGND 0.013587f
C5955 VDPWR.t540 VGND 0.013587f
C5956 VDPWR.n1390 VGND 0.029044f
C5957 VDPWR.n1391 VGND 0.11712f
C5958 VDPWR.n1392 VGND 0.116895f
C5959 VDPWR.n1393 VGND 0.028487f
C5960 VDPWR.n1394 VGND 0.175377f
C5961 VDPWR.n1395 VGND 0.078464f
C5962 VDPWR.n1396 VGND 0.052249f
C5963 VDPWR.n1397 VGND 0.158504f
C5964 VDPWR.n1398 VGND 0.052249f
C5965 VDPWR.n1399 VGND 0.207888f
C5966 VDPWR.t350 VGND 0.185586f
C5967 VDPWR.t486 VGND 0.140185f
C5968 VDPWR.t480 VGND 0.140185f
C5969 VDPWR.t352 VGND 0.186382f
C5970 VDPWR.t305 VGND 0.140185f
C5971 VDPWR.t307 VGND 0.140185f
C5972 VDPWR.t303 VGND 0.183196f
C5973 VDPWR.n1400 VGND 0.11629f
C5974 VDPWR.n1401 VGND 0.185107f
C5975 VDPWR.t518 VGND 0.186382f
C5976 VDPWR.t75 VGND 0.140185f
C5977 VDPWR.t530 VGND 0.140185f
C5978 VDPWR.t374 VGND 0.185586f
C5979 VDPWR.n1402 VGND 0.052249f
C5980 VDPWR.n1403 VGND 0.207888f
C5981 VDPWR.n1404 VGND 0.052249f
C5982 VDPWR.n1405 VGND 0.158504f
C5983 VDPWR.t120 VGND 0.185586f
C5984 VDPWR.t151 VGND 0.140185f
C5985 VDPWR.t157 VGND 0.140185f
C5986 VDPWR.t541 VGND 0.183196f
C5987 VDPWR.n1406 VGND 0.11629f
C5988 VDPWR.n1407 VGND 0.185107f
C5989 VDPWR.n1408 VGND 0.007123f
C5990 VDPWR.n1409 VGND 0.175377f
C5991 VDPWR.n1410 VGND 0.028487f
C5992 VDPWR.n1411 VGND 0.116895f
C5993 VDPWR.n1412 VGND 0.11712f
C5994 VDPWR.n1413 VGND 0.062919f
C5995 VDPWR.n1414 VGND 0.062919f
C5996 VDPWR.n1415 VGND 0.11712f
C5997 VDPWR.n1416 VGND 0.117495f
C5998 VDPWR.t304 VGND 0.013587f
C5999 VDPWR.t308 VGND 0.013587f
C6000 VDPWR.n1417 VGND 0.029044f
C6001 VDPWR.t306 VGND 0.013587f
C6002 VDPWR.t380 VGND 0.013587f
C6003 VDPWR.n1418 VGND 0.029044f
C6004 VDPWR.n1419 VGND 0.11712f
C6005 VDPWR.n1420 VGND 0.116895f
C6006 VDPWR.n1421 VGND 0.028487f
C6007 VDPWR.n1422 VGND 0.175377f
C6008 VDPWR.n1423 VGND 0.078464f
C6009 VDPWR.n1424 VGND 0.052249f
C6010 VDPWR.n1425 VGND 0.158504f
C6011 VDPWR.n1426 VGND 0.052249f
C6012 VDPWR.n1427 VGND 0.207888f
C6013 VDPWR.t584 VGND 0.185586f
C6014 VDPWR.t271 VGND 0.140185f
C6015 VDPWR.t343 VGND 0.140185f
C6016 VDPWR.t275 VGND 0.186382f
C6017 VDPWR.t89 VGND 0.140185f
C6018 VDPWR.t91 VGND 0.140185f
C6019 VDPWR.t412 VGND 0.183196f
C6020 VDPWR.n1428 VGND 0.11629f
C6021 VDPWR.n1429 VGND 0.185107f
C6022 VDPWR.t126 VGND 0.186382f
C6023 VDPWR.t73 VGND 0.140185f
C6024 VDPWR.t365 VGND 0.140185f
C6025 VDPWR.t87 VGND 0.185586f
C6026 VDPWR.n1430 VGND 0.052249f
C6027 VDPWR.n1431 VGND 0.207888f
C6028 VDPWR.n1432 VGND 0.052249f
C6029 VDPWR.n1433 VGND 0.158504f
C6030 VDPWR.t212 VGND 0.185586f
C6031 VDPWR.t313 VGND 0.140185f
C6032 VDPWR.t95 VGND 0.140185f
C6033 VDPWR.t39 VGND 0.183196f
C6034 VDPWR.n1434 VGND 0.11629f
C6035 VDPWR.n1435 VGND 0.185107f
C6036 VDPWR.n1436 VGND 0.007123f
C6037 VDPWR.n1437 VGND 0.175377f
C6038 VDPWR.n1438 VGND 0.028487f
C6039 VDPWR.n1439 VGND 0.116895f
C6040 VDPWR.n1440 VGND 0.11712f
C6041 VDPWR.n1441 VGND 0.062919f
C6042 VDPWR.n1442 VGND 0.062919f
C6043 VDPWR.n1443 VGND 0.11712f
C6044 VDPWR.n1444 VGND 0.117495f
C6045 VDPWR.t413 VGND 0.013587f
C6046 VDPWR.t92 VGND 0.013587f
C6047 VDPWR.n1445 VGND 0.029044f
C6048 VDPWR.t90 VGND 0.013587f
C6049 VDPWR.t415 VGND 0.013587f
C6050 VDPWR.n1446 VGND 0.029044f
C6051 VDPWR.n1447 VGND 0.11712f
C6052 VDPWR.n1448 VGND 0.116895f
C6053 VDPWR.n1449 VGND 0.028487f
C6054 VDPWR.n1450 VGND 0.175377f
C6055 VDPWR.n1451 VGND 0.078464f
C6056 VDPWR.n1452 VGND 0.052249f
C6057 VDPWR.n1453 VGND 0.158504f
C6058 VDPWR.n1454 VGND 0.052249f
C6059 VDPWR.n1455 VGND 0.207888f
C6060 VDPWR.t53 VGND 0.185586f
C6061 VDPWR.t422 VGND 0.140185f
C6062 VDPWR.t420 VGND 0.140185f
C6063 VDPWR.t299 VGND 0.186382f
C6064 VDPWR.n1456 VGND 0.052559f
C6065 VDPWR.n1457 VGND 0.158504f
C6066 VDPWR.t229 VGND 0.185586f
C6067 VDPWR.t200 VGND 0.140185f
C6068 VDPWR.t49 VGND 0.140185f
C6069 VDPWR.t505 VGND 0.183196f
C6070 VDPWR.n1458 VGND 0.11629f
C6071 VDPWR.n1459 VGND 0.185107f
C6072 VDPWR.n1460 VGND 0.007123f
C6073 VDPWR.n1461 VGND 0.175066f
C6074 VDPWR.n1462 VGND 0.028487f
C6075 VDPWR.n1463 VGND 0.116895f
C6076 VDPWR.n1464 VGND 0.11712f
C6077 VDPWR.n1465 VGND 0.058871f
C6078 VDPWR.n1466 VGND 0.047195f
C6079 VDPWR.t83 VGND 0.05099f
C6080 VDPWR.n1467 VGND 0.094073f
C6081 VDPWR.n1468 VGND 0.041613f
C6082 VDPWR.n1469 VGND 0.043998f
C6083 VDPWR.n1470 VGND 0.02174f
C6084 VDPWR.n1471 VGND 0.031242f
C6085 VDPWR.n1472 VGND 0.052314f
C6086 VDPWR.t198 VGND 0.05099f
C6087 VDPWR.n1473 VGND 0.043998f
C6088 VDPWR.t326 VGND 0.05099f
C6089 VDPWR.n1474 VGND 0.094073f
C6090 VDPWR.n1475 VGND 0.02174f
C6091 VDPWR.n1476 VGND 0.043998f
C6092 VDPWR.n1477 VGND 0.02174f
C6093 VDPWR.n1478 VGND 0.031242f
C6094 VDPWR.n1479 VGND 0.052314f
C6095 VDPWR.t160 VGND 0.05099f
C6096 VDPWR.n1480 VGND 0.043998f
C6097 VDPWR.t162 VGND 0.05099f
C6098 VDPWR.n1481 VGND 0.094073f
C6099 VDPWR.n1482 VGND 0.02174f
C6100 VDPWR.n1483 VGND 0.043998f
C6101 VDPWR.n1484 VGND 0.02174f
C6102 VDPWR.n1485 VGND 0.031242f
C6103 VDPWR.n1486 VGND 0.052314f
C6104 VDPWR.t159 VGND 0.05099f
C6105 VDPWR.n1487 VGND 0.010645f
C6106 VDPWR.n1488 VGND 0.031242f
C6107 VDPWR.t82 VGND 1.4182f
C6108 VDPWR.n1489 VGND 0.03114f
C6109 VDPWR.n1490 VGND 0.031242f
C6110 VDPWR.n1491 VGND 0.027943f
C6111 VDPWR.n1492 VGND 0.031242f
C6112 VDPWR.n1493 VGND 0.027943f
C6113 VDPWR.n1494 VGND 0.031242f
C6114 VDPWR.n1495 VGND 0.027943f
C6115 VDPWR.n1496 VGND 0.031242f
C6116 VDPWR.n1497 VGND 0.027943f
C6117 VDPWR.n1498 VGND 0.031242f
C6118 VDPWR.n1499 VGND 0.027943f
C6119 VDPWR.n1500 VGND 0.03114f
C6120 VDPWR.n1501 VGND 1.05038f
C6121 VDPWR.n1502 VGND 0.031242f
C6122 VDPWR.t161 VGND 0.051121f
C6123 VDPWR.n1503 VGND 0.095592f
C6124 VDPWR.n1504 VGND 0.052131f
C6125 VDPWR.n1505 VGND 0.02174f
C6126 VDPWR.n1506 VGND 0.02174f
C6127 VDPWR.n1507 VGND 0.041613f
C6128 VDPWR.n1508 VGND 0.049252f
C6129 VDPWR.n1509 VGND 0.044634f
C6130 VDPWR.t469 VGND 0.051121f
C6131 VDPWR.n1510 VGND 0.095592f
C6132 VDPWR.n1511 VGND 0.010645f
C6133 VDPWR.n1512 VGND 0.041613f
C6134 VDPWR.n1513 VGND 0.031242f
C6135 VDPWR.n1514 VGND 0.046055f
C6136 VDPWR.n1515 VGND 0.027943f
C6137 VDPWR.n1516 VGND 0.777357f
C6138 VDPWR.n1517 VGND 0.027943f
C6139 VDPWR.n1518 VGND 0.046055f
C6140 VDPWR.n1519 VGND 0.053855f
C6141 VDPWR.n1520 VGND 0.092274f
C6142 VDPWR.n1521 VGND 0.014168f
C6143 VDPWR.n1522 VGND 0.02174f
C6144 VDPWR.n1523 VGND 0.031242f
C6145 VDPWR.n1524 VGND 0.02174f
C6146 VDPWR.n1525 VGND 0.014168f
C6147 VDPWR.n1526 VGND 0.052314f
C6148 VDPWR.n1527 VGND 0.094073f
C6149 VDPWR.n1528 VGND 0.014168f
C6150 VDPWR.n1529 VGND 0.02174f
C6151 VDPWR.n1530 VGND 0.031242f
C6152 VDPWR.n1531 VGND 0.02174f
C6153 VDPWR.n1532 VGND 0.014168f
C6154 VDPWR.n1533 VGND 0.052314f
C6155 VDPWR.n1534 VGND 0.094073f
C6156 VDPWR.n1535 VGND 0.014168f
C6157 VDPWR.n1536 VGND 0.02174f
C6158 VDPWR.n1537 VGND 0.031242f
C6159 VDPWR.n1538 VGND 0.041613f
C6160 VDPWR.n1539 VGND 0.014168f
C6161 VDPWR.n1540 VGND 0.04894f
C6162 VDPWR.n1541 VGND 0.967942f
C6163 VDPWR.n1542 VGND 21.6074f
C6164 VDPWR.n1543 VGND 5.6821f
C6165 VDPWR.n1544 VGND 5.95253f
C6166 VDPWR.n1545 VGND 0.198546f
C6167 VDPWR.n1546 VGND 0.063158f
C6168 VDPWR.n1547 VGND 0.019907f
C6169 VDPWR.n1548 VGND 0.162828f
C6170 VDPWR.n1549 VGND 0.032452f
C6171 VDPWR.n1550 VGND 0.050614f
C6172 VDPWR.n1551 VGND 0.082273f
C6173 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 VGND 0.059856f
C6174 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VGND 0.019094f
C6175 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 VGND 0.041709f
C6176 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 VGND 0.059856f
C6177 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 VGND 0.019094f
C6178 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 VGND 0.04198f
C6179 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 VGND 0.013454f
C6180 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 VGND 0.059856f
C6181 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 VGND 0.019094f
C6182 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 VGND 0.04198f
C6183 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 VGND 0.059856f
C6184 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 VGND 0.019094f
C6185 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 VGND 0.041709f
C6186 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 VGND 0.013307f
C6187 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 VGND 0.351257f
C6188 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VGND 0.047903f
C6189 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 VGND 0.144997f
C6190 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 VGND 0.368007f
C6191 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 VGND 0.013091f
C6192 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 VGND 0.013091f
C6193 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 VGND 0.030662f
C6194 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 VGND 0.039272f
C6195 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 VGND 0.039272f
C6196 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 VGND 0.080004f
C6197 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 VGND 0.332866f
C6198 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 VGND 0.060722f
C6199 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 VGND 0.060722f
C6200 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 VGND 0.070899f
C6201 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 VGND 0.060722f
C6202 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 VGND 0.060722f
C6203 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 VGND 0.070523f
C6204 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 VGND 0.632153f
C6205 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 VGND 0.045973f
C6206 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 VGND 0.156775f
C6207 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 VGND 0.144997f
C6208 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 VGND 0.240639f
C6209 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 VGND 0.180864f
.ends

