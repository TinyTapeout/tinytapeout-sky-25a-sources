magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -415 -300 415 300
<< nmos >>
rect -229 -100 -29 100
rect 29 -100 229 100
<< ndiff >>
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
<< ndiffc >>
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
<< psubdiff >>
rect -389 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 389 274
rect -389 153 -355 240
rect -389 85 -355 119
rect 355 153 389 240
rect -389 17 -355 51
rect -389 -51 -355 -17
rect -389 -119 -355 -85
rect 355 85 389 119
rect 355 17 389 51
rect 355 -51 389 -17
rect -389 -240 -355 -153
rect 355 -119 389 -85
rect 355 -240 389 -153
rect -389 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 389 -240
<< psubdiffcont >>
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect -389 119 -355 153
rect 355 119 389 153
rect -389 51 -355 85
rect -389 -17 -355 17
rect -389 -85 -355 -51
rect 355 51 389 85
rect 355 -17 389 17
rect 355 -85 389 -51
rect -389 -153 -355 -119
rect 355 -153 389 -119
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
<< poly >>
rect -229 172 -29 188
rect -229 138 -180 172
rect -146 138 -112 172
rect -78 138 -29 172
rect -229 100 -29 138
rect 29 172 229 188
rect 29 138 78 172
rect 112 138 146 172
rect 180 138 229 172
rect 29 100 229 138
rect -229 -138 -29 -100
rect -229 -172 -180 -138
rect -146 -172 -112 -138
rect -78 -172 -29 -138
rect -229 -188 -29 -172
rect 29 -138 229 -100
rect 29 -172 78 -138
rect 112 -172 146 -138
rect 180 -172 229 -138
rect 29 -188 229 -172
<< polycont >>
rect -180 138 -146 172
rect -112 138 -78 172
rect 78 138 112 172
rect 146 138 180 172
rect -180 -172 -146 -138
rect -112 -172 -78 -138
rect 78 -172 112 -138
rect 146 -172 180 -138
<< locali >>
rect -389 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 389 274
rect -389 153 -355 240
rect -229 138 -182 172
rect -146 138 -112 172
rect -76 138 -29 172
rect 29 138 76 172
rect 112 138 146 172
rect 182 138 229 172
rect 355 153 389 240
rect -389 85 -355 119
rect -389 17 -355 51
rect -389 -51 -355 -17
rect -389 -119 -355 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 355 85 389 119
rect 355 17 389 51
rect 355 -51 389 -17
rect 355 -119 389 -85
rect -389 -240 -355 -153
rect -229 -172 -182 -138
rect -146 -172 -112 -138
rect -76 -172 -29 -138
rect 29 -172 76 -138
rect 112 -172 146 -138
rect 182 -172 229 -138
rect 355 -240 389 -153
rect -389 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 389 -240
<< viali >>
rect -182 138 -180 172
rect -180 138 -148 172
rect -110 138 -78 172
rect -78 138 -76 172
rect 76 138 78 172
rect 78 138 110 172
rect 148 138 180 172
rect 180 138 182 172
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect -182 -172 -180 -138
rect -180 -172 -148 -138
rect -110 -172 -78 -138
rect -78 -172 -76 -138
rect 76 -172 78 -138
rect 78 -172 110 -138
rect 148 -172 180 -138
rect 180 -172 182 -138
<< metal1 >>
rect -225 172 -33 178
rect -225 138 -182 172
rect -148 138 -110 172
rect -76 138 -33 172
rect -225 132 -33 138
rect 33 172 225 178
rect 33 138 76 172
rect 110 138 148 172
rect 182 138 225 172
rect 33 132 225 138
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect -225 -138 -33 -132
rect -225 -172 -182 -138
rect -148 -172 -110 -138
rect -76 -172 -33 -138
rect -225 -178 -33 -172
rect 33 -138 225 -132
rect 33 -172 76 -138
rect 110 -172 148 -138
rect 182 -172 225 -138
rect 33 -178 225 -172
<< properties >>
string FIXED_BBOX -372 -257 372 257
<< end >>
