magic
tech sky130A
magscale 1 2
timestamp 1757256469
<< pwell >>
rect -1781 -327 1781 327
<< mvnmos >>
rect -1551 -131 -1451 69
rect -1393 -131 -1293 69
rect -1235 -131 -1135 69
rect -1077 -131 -977 69
rect -919 -131 -819 69
rect -761 -131 -661 69
rect -603 -131 -503 69
rect -445 -131 -345 69
rect -287 -131 -187 69
rect -129 -131 -29 69
rect 29 -131 129 69
rect 187 -131 287 69
rect 345 -131 445 69
rect 503 -131 603 69
rect 661 -131 761 69
rect 819 -131 919 69
rect 977 -131 1077 69
rect 1135 -131 1235 69
rect 1293 -131 1393 69
rect 1451 -131 1551 69
<< mvndiff >>
rect -1609 57 -1551 69
rect -1609 -119 -1597 57
rect -1563 -119 -1551 57
rect -1609 -131 -1551 -119
rect -1451 57 -1393 69
rect -1451 -119 -1439 57
rect -1405 -119 -1393 57
rect -1451 -131 -1393 -119
rect -1293 57 -1235 69
rect -1293 -119 -1281 57
rect -1247 -119 -1235 57
rect -1293 -131 -1235 -119
rect -1135 57 -1077 69
rect -1135 -119 -1123 57
rect -1089 -119 -1077 57
rect -1135 -131 -1077 -119
rect -977 57 -919 69
rect -977 -119 -965 57
rect -931 -119 -919 57
rect -977 -131 -919 -119
rect -819 57 -761 69
rect -819 -119 -807 57
rect -773 -119 -761 57
rect -819 -131 -761 -119
rect -661 57 -603 69
rect -661 -119 -649 57
rect -615 -119 -603 57
rect -661 -131 -603 -119
rect -503 57 -445 69
rect -503 -119 -491 57
rect -457 -119 -445 57
rect -503 -131 -445 -119
rect -345 57 -287 69
rect -345 -119 -333 57
rect -299 -119 -287 57
rect -345 -131 -287 -119
rect -187 57 -129 69
rect -187 -119 -175 57
rect -141 -119 -129 57
rect -187 -131 -129 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 129 57 187 69
rect 129 -119 141 57
rect 175 -119 187 57
rect 129 -131 187 -119
rect 287 57 345 69
rect 287 -119 299 57
rect 333 -119 345 57
rect 287 -131 345 -119
rect 445 57 503 69
rect 445 -119 457 57
rect 491 -119 503 57
rect 445 -131 503 -119
rect 603 57 661 69
rect 603 -119 615 57
rect 649 -119 661 57
rect 603 -131 661 -119
rect 761 57 819 69
rect 761 -119 773 57
rect 807 -119 819 57
rect 761 -131 819 -119
rect 919 57 977 69
rect 919 -119 931 57
rect 965 -119 977 57
rect 919 -131 977 -119
rect 1077 57 1135 69
rect 1077 -119 1089 57
rect 1123 -119 1135 57
rect 1077 -131 1135 -119
rect 1235 57 1293 69
rect 1235 -119 1247 57
rect 1281 -119 1293 57
rect 1235 -131 1293 -119
rect 1393 57 1451 69
rect 1393 -119 1405 57
rect 1439 -119 1451 57
rect 1393 -131 1451 -119
rect 1551 57 1609 69
rect 1551 -119 1563 57
rect 1597 -119 1609 57
rect 1551 -131 1609 -119
<< mvndiffc >>
rect -1597 -119 -1563 57
rect -1439 -119 -1405 57
rect -1281 -119 -1247 57
rect -1123 -119 -1089 57
rect -965 -119 -931 57
rect -807 -119 -773 57
rect -649 -119 -615 57
rect -491 -119 -457 57
rect -333 -119 -299 57
rect -175 -119 -141 57
rect -17 -119 17 57
rect 141 -119 175 57
rect 299 -119 333 57
rect 457 -119 491 57
rect 615 -119 649 57
rect 773 -119 807 57
rect 931 -119 965 57
rect 1089 -119 1123 57
rect 1247 -119 1281 57
rect 1405 -119 1439 57
rect 1563 -119 1597 57
<< mvpsubdiff >>
rect -1745 279 1745 291
rect -1745 245 -1637 279
rect 1637 245 1745 279
rect -1745 233 1745 245
rect -1745 183 -1687 233
rect -1745 -183 -1733 183
rect -1699 -183 -1687 183
rect 1687 183 1745 233
rect -1745 -233 -1687 -183
rect 1687 -183 1699 183
rect 1733 -183 1745 183
rect 1687 -233 1745 -183
rect -1745 -245 1745 -233
rect -1745 -279 -1637 -245
rect 1637 -279 1745 -245
rect -1745 -291 1745 -279
<< mvpsubdiffcont >>
rect -1637 245 1637 279
rect -1733 -183 -1699 183
rect 1699 -183 1733 183
rect -1637 -279 1637 -245
<< poly >>
rect -1551 141 -1451 157
rect -1551 107 -1535 141
rect -1467 107 -1451 141
rect -1551 69 -1451 107
rect -1393 141 -1293 157
rect -1393 107 -1377 141
rect -1309 107 -1293 141
rect -1393 69 -1293 107
rect -1235 141 -1135 157
rect -1235 107 -1219 141
rect -1151 107 -1135 141
rect -1235 69 -1135 107
rect -1077 141 -977 157
rect -1077 107 -1061 141
rect -993 107 -977 141
rect -1077 69 -977 107
rect -919 141 -819 157
rect -919 107 -903 141
rect -835 107 -819 141
rect -919 69 -819 107
rect -761 141 -661 157
rect -761 107 -745 141
rect -677 107 -661 141
rect -761 69 -661 107
rect -603 141 -503 157
rect -603 107 -587 141
rect -519 107 -503 141
rect -603 69 -503 107
rect -445 141 -345 157
rect -445 107 -429 141
rect -361 107 -345 141
rect -445 69 -345 107
rect -287 141 -187 157
rect -287 107 -271 141
rect -203 107 -187 141
rect -287 69 -187 107
rect -129 141 -29 157
rect -129 107 -113 141
rect -45 107 -29 141
rect -129 69 -29 107
rect 29 141 129 157
rect 29 107 45 141
rect 113 107 129 141
rect 29 69 129 107
rect 187 141 287 157
rect 187 107 203 141
rect 271 107 287 141
rect 187 69 287 107
rect 345 141 445 157
rect 345 107 361 141
rect 429 107 445 141
rect 345 69 445 107
rect 503 141 603 157
rect 503 107 519 141
rect 587 107 603 141
rect 503 69 603 107
rect 661 141 761 157
rect 661 107 677 141
rect 745 107 761 141
rect 661 69 761 107
rect 819 141 919 157
rect 819 107 835 141
rect 903 107 919 141
rect 819 69 919 107
rect 977 141 1077 157
rect 977 107 993 141
rect 1061 107 1077 141
rect 977 69 1077 107
rect 1135 141 1235 157
rect 1135 107 1151 141
rect 1219 107 1235 141
rect 1135 69 1235 107
rect 1293 141 1393 157
rect 1293 107 1309 141
rect 1377 107 1393 141
rect 1293 69 1393 107
rect 1451 141 1551 157
rect 1451 107 1467 141
rect 1535 107 1551 141
rect 1451 69 1551 107
rect -1551 -157 -1451 -131
rect -1393 -157 -1293 -131
rect -1235 -157 -1135 -131
rect -1077 -157 -977 -131
rect -919 -157 -819 -131
rect -761 -157 -661 -131
rect -603 -157 -503 -131
rect -445 -157 -345 -131
rect -287 -157 -187 -131
rect -129 -157 -29 -131
rect 29 -157 129 -131
rect 187 -157 287 -131
rect 345 -157 445 -131
rect 503 -157 603 -131
rect 661 -157 761 -131
rect 819 -157 919 -131
rect 977 -157 1077 -131
rect 1135 -157 1235 -131
rect 1293 -157 1393 -131
rect 1451 -157 1551 -131
<< polycont >>
rect -1535 107 -1467 141
rect -1377 107 -1309 141
rect -1219 107 -1151 141
rect -1061 107 -993 141
rect -903 107 -835 141
rect -745 107 -677 141
rect -587 107 -519 141
rect -429 107 -361 141
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
rect 361 107 429 141
rect 519 107 587 141
rect 677 107 745 141
rect 835 107 903 141
rect 993 107 1061 141
rect 1151 107 1219 141
rect 1309 107 1377 141
rect 1467 107 1535 141
<< locali >>
rect -1733 245 -1637 279
rect 1637 245 1733 279
rect -1733 183 -1699 245
rect 1699 183 1733 245
rect -1551 107 -1535 141
rect -1467 107 -1451 141
rect -1393 107 -1377 141
rect -1309 107 -1293 141
rect -1235 107 -1219 141
rect -1151 107 -1135 141
rect -1077 107 -1061 141
rect -993 107 -977 141
rect -919 107 -903 141
rect -835 107 -819 141
rect -761 107 -745 141
rect -677 107 -661 141
rect -603 107 -587 141
rect -519 107 -503 141
rect -445 107 -429 141
rect -361 107 -345 141
rect -287 107 -271 141
rect -203 107 -187 141
rect -129 107 -113 141
rect -45 107 -29 141
rect 29 107 45 141
rect 113 107 129 141
rect 187 107 203 141
rect 271 107 287 141
rect 345 107 361 141
rect 429 107 445 141
rect 503 107 519 141
rect 587 107 603 141
rect 661 107 677 141
rect 745 107 761 141
rect 819 107 835 141
rect 903 107 919 141
rect 977 107 993 141
rect 1061 107 1077 141
rect 1135 107 1151 141
rect 1219 107 1235 141
rect 1293 107 1309 141
rect 1377 107 1393 141
rect 1451 107 1467 141
rect 1535 107 1551 141
rect -1597 57 -1563 73
rect -1597 -135 -1563 -119
rect -1439 57 -1405 73
rect -1439 -135 -1405 -119
rect -1281 57 -1247 73
rect -1281 -135 -1247 -119
rect -1123 57 -1089 73
rect -1123 -135 -1089 -119
rect -965 57 -931 73
rect -965 -135 -931 -119
rect -807 57 -773 73
rect -807 -135 -773 -119
rect -649 57 -615 73
rect -649 -135 -615 -119
rect -491 57 -457 73
rect -491 -135 -457 -119
rect -333 57 -299 73
rect -333 -135 -299 -119
rect -175 57 -141 73
rect -175 -135 -141 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 141 57 175 73
rect 141 -135 175 -119
rect 299 57 333 73
rect 299 -135 333 -119
rect 457 57 491 73
rect 457 -135 491 -119
rect 615 57 649 73
rect 615 -135 649 -119
rect 773 57 807 73
rect 773 -135 807 -119
rect 931 57 965 73
rect 931 -135 965 -119
rect 1089 57 1123 73
rect 1089 -135 1123 -119
rect 1247 57 1281 73
rect 1247 -135 1281 -119
rect 1405 57 1439 73
rect 1405 -135 1439 -119
rect 1563 57 1597 73
rect 1563 -135 1597 -119
rect -1733 -245 -1699 -183
rect 1699 -245 1733 -183
rect -1733 -279 -1637 -245
rect 1637 -279 1733 -245
<< viali >>
rect -1535 107 -1467 141
rect -1377 107 -1309 141
rect -1219 107 -1151 141
rect -1061 107 -993 141
rect -903 107 -835 141
rect -745 107 -677 141
rect -587 107 -519 141
rect -429 107 -361 141
rect -271 107 -203 141
rect -113 107 -45 141
rect 45 107 113 141
rect 203 107 271 141
rect 361 107 429 141
rect 519 107 587 141
rect 677 107 745 141
rect 835 107 903 141
rect 993 107 1061 141
rect 1151 107 1219 141
rect 1309 107 1377 141
rect 1467 107 1535 141
rect -1597 -119 -1563 57
rect -1439 -119 -1405 57
rect -1281 -119 -1247 57
rect -1123 -119 -1089 57
rect -965 -119 -931 57
rect -807 -119 -773 57
rect -649 -119 -615 57
rect -491 -119 -457 57
rect -333 -119 -299 57
rect -175 -119 -141 57
rect -17 -119 17 57
rect 141 -119 175 57
rect 299 -119 333 57
rect 457 -119 491 57
rect 615 -119 649 57
rect 773 -119 807 57
rect 931 -119 965 57
rect 1089 -119 1123 57
rect 1247 -119 1281 57
rect 1405 -119 1439 57
rect 1563 -119 1597 57
<< metal1 >>
rect -1547 141 -1455 147
rect -1547 107 -1535 141
rect -1467 107 -1455 141
rect -1547 101 -1455 107
rect -1389 141 -1297 147
rect -1389 107 -1377 141
rect -1309 107 -1297 141
rect -1389 101 -1297 107
rect -1231 141 -1139 147
rect -1231 107 -1219 141
rect -1151 107 -1139 141
rect -1231 101 -1139 107
rect -1073 141 -981 147
rect -1073 107 -1061 141
rect -993 107 -981 141
rect -1073 101 -981 107
rect -915 141 -823 147
rect -915 107 -903 141
rect -835 107 -823 141
rect -915 101 -823 107
rect -757 141 -665 147
rect -757 107 -745 141
rect -677 107 -665 141
rect -757 101 -665 107
rect -599 141 -507 147
rect -599 107 -587 141
rect -519 107 -507 141
rect -599 101 -507 107
rect -441 141 -349 147
rect -441 107 -429 141
rect -361 107 -349 141
rect -441 101 -349 107
rect -283 141 -191 147
rect -283 107 -271 141
rect -203 107 -191 141
rect -283 101 -191 107
rect -125 141 -33 147
rect -125 107 -113 141
rect -45 107 -33 141
rect -125 101 -33 107
rect 33 141 125 147
rect 33 107 45 141
rect 113 107 125 141
rect 33 101 125 107
rect 191 141 283 147
rect 191 107 203 141
rect 271 107 283 141
rect 191 101 283 107
rect 349 141 441 147
rect 349 107 361 141
rect 429 107 441 141
rect 349 101 441 107
rect 507 141 599 147
rect 507 107 519 141
rect 587 107 599 141
rect 507 101 599 107
rect 665 141 757 147
rect 665 107 677 141
rect 745 107 757 141
rect 665 101 757 107
rect 823 141 915 147
rect 823 107 835 141
rect 903 107 915 141
rect 823 101 915 107
rect 981 141 1073 147
rect 981 107 993 141
rect 1061 107 1073 141
rect 981 101 1073 107
rect 1139 141 1231 147
rect 1139 107 1151 141
rect 1219 107 1231 141
rect 1139 101 1231 107
rect 1297 141 1389 147
rect 1297 107 1309 141
rect 1377 107 1389 141
rect 1297 101 1389 107
rect 1455 141 1547 147
rect 1455 107 1467 141
rect 1535 107 1547 141
rect 1455 101 1547 107
rect -1603 57 -1557 69
rect -1603 -119 -1597 57
rect -1563 -119 -1557 57
rect -1603 -131 -1557 -119
rect -1445 57 -1399 69
rect -1445 -119 -1439 57
rect -1405 -119 -1399 57
rect -1445 -131 -1399 -119
rect -1287 57 -1241 69
rect -1287 -119 -1281 57
rect -1247 -119 -1241 57
rect -1287 -131 -1241 -119
rect -1129 57 -1083 69
rect -1129 -119 -1123 57
rect -1089 -119 -1083 57
rect -1129 -131 -1083 -119
rect -971 57 -925 69
rect -971 -119 -965 57
rect -931 -119 -925 57
rect -971 -131 -925 -119
rect -813 57 -767 69
rect -813 -119 -807 57
rect -773 -119 -767 57
rect -813 -131 -767 -119
rect -655 57 -609 69
rect -655 -119 -649 57
rect -615 -119 -609 57
rect -655 -131 -609 -119
rect -497 57 -451 69
rect -497 -119 -491 57
rect -457 -119 -451 57
rect -497 -131 -451 -119
rect -339 57 -293 69
rect -339 -119 -333 57
rect -299 -119 -293 57
rect -339 -131 -293 -119
rect -181 57 -135 69
rect -181 -119 -175 57
rect -141 -119 -135 57
rect -181 -131 -135 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 135 57 181 69
rect 135 -119 141 57
rect 175 -119 181 57
rect 135 -131 181 -119
rect 293 57 339 69
rect 293 -119 299 57
rect 333 -119 339 57
rect 293 -131 339 -119
rect 451 57 497 69
rect 451 -119 457 57
rect 491 -119 497 57
rect 451 -131 497 -119
rect 609 57 655 69
rect 609 -119 615 57
rect 649 -119 655 57
rect 609 -131 655 -119
rect 767 57 813 69
rect 767 -119 773 57
rect 807 -119 813 57
rect 767 -131 813 -119
rect 925 57 971 69
rect 925 -119 931 57
rect 965 -119 971 57
rect 925 -131 971 -119
rect 1083 57 1129 69
rect 1083 -119 1089 57
rect 1123 -119 1129 57
rect 1083 -131 1129 -119
rect 1241 57 1287 69
rect 1241 -119 1247 57
rect 1281 -119 1287 57
rect 1241 -131 1287 -119
rect 1399 57 1445 69
rect 1399 -119 1405 57
rect 1439 -119 1445 57
rect 1399 -131 1445 -119
rect 1557 57 1603 69
rect 1557 -119 1563 57
rect 1597 -119 1603 57
rect 1557 -131 1603 -119
<< labels >>
rlabel mvpsubdiffcont 0 -262 0 -262 0 B
port 1 nsew
rlabel mvndiffc -1580 -31 -1580 -31 0 D0
port 2 nsew
rlabel polycont -1501 124 -1501 124 0 G0
port 3 nsew
rlabel mvndiffc -1422 -31 -1422 -31 0 S1
port 4 nsew
rlabel polycont -1343 124 -1343 124 0 G1
port 5 nsew
rlabel mvndiffc -1264 -31 -1264 -31 0 D2
port 6 nsew
rlabel polycont -1185 124 -1185 124 0 G2
port 7 nsew
rlabel mvndiffc -1106 -31 -1106 -31 0 S3
port 8 nsew
rlabel polycont -1027 124 -1027 124 0 G3
port 9 nsew
rlabel mvndiffc -948 -31 -948 -31 0 D4
port 10 nsew
rlabel polycont -869 124 -869 124 0 G4
port 11 nsew
rlabel mvndiffc -790 -31 -790 -31 0 S5
port 12 nsew
rlabel polycont -711 124 -711 124 0 G5
port 13 nsew
rlabel mvndiffc -632 -31 -632 -31 0 D6
port 14 nsew
rlabel polycont -553 124 -553 124 0 G6
port 15 nsew
rlabel mvndiffc -474 -31 -474 -31 0 S7
port 16 nsew
rlabel polycont -395 124 -395 124 0 G7
port 17 nsew
rlabel mvndiffc -316 -31 -316 -31 0 D8
port 18 nsew
rlabel polycont -237 124 -237 124 0 G8
port 19 nsew
rlabel mvndiffc -158 -31 -158 -31 0 S9
port 20 nsew
rlabel polycont -79 124 -79 124 0 G9
port 21 nsew
rlabel mvndiffc 0 -31 0 -31 0 D10
port 22 nsew
rlabel polycont 79 124 79 124 0 G10
port 23 nsew
rlabel mvndiffc 158 -31 158 -31 0 S11
port 24 nsew
rlabel polycont 237 124 237 124 0 G11
port 25 nsew
rlabel mvndiffc 316 -31 316 -31 0 D12
port 26 nsew
rlabel polycont 395 124 395 124 0 G12
port 27 nsew
rlabel mvndiffc 474 -31 474 -31 0 S13
port 28 nsew
rlabel polycont 553 124 553 124 0 G13
port 29 nsew
rlabel mvndiffc 632 -31 632 -31 0 D14
port 30 nsew
rlabel polycont 711 124 711 124 0 G14
port 31 nsew
rlabel mvndiffc 790 -31 790 -31 0 S15
port 32 nsew
rlabel polycont 869 124 869 124 0 G15
port 33 nsew
rlabel mvndiffc 948 -31 948 -31 0 D16
port 34 nsew
rlabel polycont 1027 124 1027 124 0 G16
port 35 nsew
rlabel mvndiffc 1106 -31 1106 -31 0 S17
port 36 nsew
rlabel polycont 1185 124 1185 124 0 G17
port 37 nsew
rlabel mvndiffc 1264 -31 1264 -31 0 D18
port 38 nsew
rlabel polycont 1343 124 1343 124 0 G18
port 39 nsew
rlabel mvndiffc 1422 -31 1422 -31 0 S19
port 40 nsew
rlabel polycont 1501 124 1501 124 0 G19
port 41 nsew
<< properties >>
string FIXED_BBOX -1716 -262 1716 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
