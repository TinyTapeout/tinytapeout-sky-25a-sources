
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* Increment toggling
Vinc INC_IN VGND pulse(0 1.8 1.5n 200p 200p 2n 4n)
Rinc INC_IN INC 100

* create clock
Vclk CLK_IN VGND pulse(0 1.8 1n 200p 200p 1n 2n)
Vrstn RSTN VGND pulse(1.8 0 100n 50p 50p 5n)
.tran 10e-12 500e-09 0e-00

Rclk CLK_IN CLK 100

Rs0 S0 S0_OUT 100
Rs1 S1 S1_OUT 100
Rs2 S2 S2_OUT 100
Rs3 S3 S3_OUT 100
Rs4 S4 S4_OUT 100
Rs5 S5 S5_OUT 100

Cs0 S0_OUT VGND 1f
Cs1 S1_OUT VGND 1f
Cs2 S2_OUT VGND 1f
Cs3 S3_OUT VGND 1f
Cs4 S4_OUT VGND 1f
Cs5 S5_OUT VGND 1f

.control
run
set color0 = white
set color1 = black
plot INC-0.4 CLK-0.2 S0_OUT S1_OUT+0.2 S2_OUT+0.4 S3_OUT+0.6 S4_OUT+0.8
plot RSTN-0.4 S0 S5+0.2 S6+0.4 S7+0.6 S8+0.8 S9+1.0
plot i(Vdd)
.endc

.end
