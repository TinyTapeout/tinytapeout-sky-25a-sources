magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -673 -1200 673 1200
<< nmos >>
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
<< ndiff >>
rect -545 969 -487 1000
rect -545 935 -533 969
rect -499 935 -487 969
rect -545 901 -487 935
rect -545 867 -533 901
rect -499 867 -487 901
rect -545 833 -487 867
rect -545 799 -533 833
rect -499 799 -487 833
rect -545 765 -487 799
rect -545 731 -533 765
rect -499 731 -487 765
rect -545 697 -487 731
rect -545 663 -533 697
rect -499 663 -487 697
rect -545 629 -487 663
rect -545 595 -533 629
rect -499 595 -487 629
rect -545 561 -487 595
rect -545 527 -533 561
rect -499 527 -487 561
rect -545 493 -487 527
rect -545 459 -533 493
rect -499 459 -487 493
rect -545 425 -487 459
rect -545 391 -533 425
rect -499 391 -487 425
rect -545 357 -487 391
rect -545 323 -533 357
rect -499 323 -487 357
rect -545 289 -487 323
rect -545 255 -533 289
rect -499 255 -487 289
rect -545 221 -487 255
rect -545 187 -533 221
rect -499 187 -487 221
rect -545 153 -487 187
rect -545 119 -533 153
rect -499 119 -487 153
rect -545 85 -487 119
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -119 -487 -85
rect -545 -153 -533 -119
rect -499 -153 -487 -119
rect -545 -187 -487 -153
rect -545 -221 -533 -187
rect -499 -221 -487 -187
rect -545 -255 -487 -221
rect -545 -289 -533 -255
rect -499 -289 -487 -255
rect -545 -323 -487 -289
rect -545 -357 -533 -323
rect -499 -357 -487 -323
rect -545 -391 -487 -357
rect -545 -425 -533 -391
rect -499 -425 -487 -391
rect -545 -459 -487 -425
rect -545 -493 -533 -459
rect -499 -493 -487 -459
rect -545 -527 -487 -493
rect -545 -561 -533 -527
rect -499 -561 -487 -527
rect -545 -595 -487 -561
rect -545 -629 -533 -595
rect -499 -629 -487 -595
rect -545 -663 -487 -629
rect -545 -697 -533 -663
rect -499 -697 -487 -663
rect -545 -731 -487 -697
rect -545 -765 -533 -731
rect -499 -765 -487 -731
rect -545 -799 -487 -765
rect -545 -833 -533 -799
rect -499 -833 -487 -799
rect -545 -867 -487 -833
rect -545 -901 -533 -867
rect -499 -901 -487 -867
rect -545 -935 -487 -901
rect -545 -969 -533 -935
rect -499 -969 -487 -935
rect -545 -1000 -487 -969
rect -287 969 -229 1000
rect -287 935 -275 969
rect -241 935 -229 969
rect -287 901 -229 935
rect -287 867 -275 901
rect -241 867 -229 901
rect -287 833 -229 867
rect -287 799 -275 833
rect -241 799 -229 833
rect -287 765 -229 799
rect -287 731 -275 765
rect -241 731 -229 765
rect -287 697 -229 731
rect -287 663 -275 697
rect -241 663 -229 697
rect -287 629 -229 663
rect -287 595 -275 629
rect -241 595 -229 629
rect -287 561 -229 595
rect -287 527 -275 561
rect -241 527 -229 561
rect -287 493 -229 527
rect -287 459 -275 493
rect -241 459 -229 493
rect -287 425 -229 459
rect -287 391 -275 425
rect -241 391 -229 425
rect -287 357 -229 391
rect -287 323 -275 357
rect -241 323 -229 357
rect -287 289 -229 323
rect -287 255 -275 289
rect -241 255 -229 289
rect -287 221 -229 255
rect -287 187 -275 221
rect -241 187 -229 221
rect -287 153 -229 187
rect -287 119 -275 153
rect -241 119 -229 153
rect -287 85 -229 119
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -119 -229 -85
rect -287 -153 -275 -119
rect -241 -153 -229 -119
rect -287 -187 -229 -153
rect -287 -221 -275 -187
rect -241 -221 -229 -187
rect -287 -255 -229 -221
rect -287 -289 -275 -255
rect -241 -289 -229 -255
rect -287 -323 -229 -289
rect -287 -357 -275 -323
rect -241 -357 -229 -323
rect -287 -391 -229 -357
rect -287 -425 -275 -391
rect -241 -425 -229 -391
rect -287 -459 -229 -425
rect -287 -493 -275 -459
rect -241 -493 -229 -459
rect -287 -527 -229 -493
rect -287 -561 -275 -527
rect -241 -561 -229 -527
rect -287 -595 -229 -561
rect -287 -629 -275 -595
rect -241 -629 -229 -595
rect -287 -663 -229 -629
rect -287 -697 -275 -663
rect -241 -697 -229 -663
rect -287 -731 -229 -697
rect -287 -765 -275 -731
rect -241 -765 -229 -731
rect -287 -799 -229 -765
rect -287 -833 -275 -799
rect -241 -833 -229 -799
rect -287 -867 -229 -833
rect -287 -901 -275 -867
rect -241 -901 -229 -867
rect -287 -935 -229 -901
rect -287 -969 -275 -935
rect -241 -969 -229 -935
rect -287 -1000 -229 -969
rect -29 969 29 1000
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1000 29 -969
rect 229 969 287 1000
rect 229 935 241 969
rect 275 935 287 969
rect 229 901 287 935
rect 229 867 241 901
rect 275 867 287 901
rect 229 833 287 867
rect 229 799 241 833
rect 275 799 287 833
rect 229 765 287 799
rect 229 731 241 765
rect 275 731 287 765
rect 229 697 287 731
rect 229 663 241 697
rect 275 663 287 697
rect 229 629 287 663
rect 229 595 241 629
rect 275 595 287 629
rect 229 561 287 595
rect 229 527 241 561
rect 275 527 287 561
rect 229 493 287 527
rect 229 459 241 493
rect 275 459 287 493
rect 229 425 287 459
rect 229 391 241 425
rect 275 391 287 425
rect 229 357 287 391
rect 229 323 241 357
rect 275 323 287 357
rect 229 289 287 323
rect 229 255 241 289
rect 275 255 287 289
rect 229 221 287 255
rect 229 187 241 221
rect 275 187 287 221
rect 229 153 287 187
rect 229 119 241 153
rect 275 119 287 153
rect 229 85 287 119
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -119 287 -85
rect 229 -153 241 -119
rect 275 -153 287 -119
rect 229 -187 287 -153
rect 229 -221 241 -187
rect 275 -221 287 -187
rect 229 -255 287 -221
rect 229 -289 241 -255
rect 275 -289 287 -255
rect 229 -323 287 -289
rect 229 -357 241 -323
rect 275 -357 287 -323
rect 229 -391 287 -357
rect 229 -425 241 -391
rect 275 -425 287 -391
rect 229 -459 287 -425
rect 229 -493 241 -459
rect 275 -493 287 -459
rect 229 -527 287 -493
rect 229 -561 241 -527
rect 275 -561 287 -527
rect 229 -595 287 -561
rect 229 -629 241 -595
rect 275 -629 287 -595
rect 229 -663 287 -629
rect 229 -697 241 -663
rect 275 -697 287 -663
rect 229 -731 287 -697
rect 229 -765 241 -731
rect 275 -765 287 -731
rect 229 -799 287 -765
rect 229 -833 241 -799
rect 275 -833 287 -799
rect 229 -867 287 -833
rect 229 -901 241 -867
rect 275 -901 287 -867
rect 229 -935 287 -901
rect 229 -969 241 -935
rect 275 -969 287 -935
rect 229 -1000 287 -969
rect 487 969 545 1000
rect 487 935 499 969
rect 533 935 545 969
rect 487 901 545 935
rect 487 867 499 901
rect 533 867 545 901
rect 487 833 545 867
rect 487 799 499 833
rect 533 799 545 833
rect 487 765 545 799
rect 487 731 499 765
rect 533 731 545 765
rect 487 697 545 731
rect 487 663 499 697
rect 533 663 545 697
rect 487 629 545 663
rect 487 595 499 629
rect 533 595 545 629
rect 487 561 545 595
rect 487 527 499 561
rect 533 527 545 561
rect 487 493 545 527
rect 487 459 499 493
rect 533 459 545 493
rect 487 425 545 459
rect 487 391 499 425
rect 533 391 545 425
rect 487 357 545 391
rect 487 323 499 357
rect 533 323 545 357
rect 487 289 545 323
rect 487 255 499 289
rect 533 255 545 289
rect 487 221 545 255
rect 487 187 499 221
rect 533 187 545 221
rect 487 153 545 187
rect 487 119 499 153
rect 533 119 545 153
rect 487 85 545 119
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -119 545 -85
rect 487 -153 499 -119
rect 533 -153 545 -119
rect 487 -187 545 -153
rect 487 -221 499 -187
rect 533 -221 545 -187
rect 487 -255 545 -221
rect 487 -289 499 -255
rect 533 -289 545 -255
rect 487 -323 545 -289
rect 487 -357 499 -323
rect 533 -357 545 -323
rect 487 -391 545 -357
rect 487 -425 499 -391
rect 533 -425 545 -391
rect 487 -459 545 -425
rect 487 -493 499 -459
rect 533 -493 545 -459
rect 487 -527 545 -493
rect 487 -561 499 -527
rect 533 -561 545 -527
rect 487 -595 545 -561
rect 487 -629 499 -595
rect 533 -629 545 -595
rect 487 -663 545 -629
rect 487 -697 499 -663
rect 533 -697 545 -663
rect 487 -731 545 -697
rect 487 -765 499 -731
rect 533 -765 545 -731
rect 487 -799 545 -765
rect 487 -833 499 -799
rect 533 -833 545 -799
rect 487 -867 545 -833
rect 487 -901 499 -867
rect 533 -901 545 -867
rect 487 -935 545 -901
rect 487 -969 499 -935
rect 533 -969 545 -935
rect 487 -1000 545 -969
<< ndiffc >>
rect -533 935 -499 969
rect -533 867 -499 901
rect -533 799 -499 833
rect -533 731 -499 765
rect -533 663 -499 697
rect -533 595 -499 629
rect -533 527 -499 561
rect -533 459 -499 493
rect -533 391 -499 425
rect -533 323 -499 357
rect -533 255 -499 289
rect -533 187 -499 221
rect -533 119 -499 153
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -533 -153 -499 -119
rect -533 -221 -499 -187
rect -533 -289 -499 -255
rect -533 -357 -499 -323
rect -533 -425 -499 -391
rect -533 -493 -499 -459
rect -533 -561 -499 -527
rect -533 -629 -499 -595
rect -533 -697 -499 -663
rect -533 -765 -499 -731
rect -533 -833 -499 -799
rect -533 -901 -499 -867
rect -533 -969 -499 -935
rect -275 935 -241 969
rect -275 867 -241 901
rect -275 799 -241 833
rect -275 731 -241 765
rect -275 663 -241 697
rect -275 595 -241 629
rect -275 527 -241 561
rect -275 459 -241 493
rect -275 391 -241 425
rect -275 323 -241 357
rect -275 255 -241 289
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -275 -289 -241 -255
rect -275 -357 -241 -323
rect -275 -425 -241 -391
rect -275 -493 -241 -459
rect -275 -561 -241 -527
rect -275 -629 -241 -595
rect -275 -697 -241 -663
rect -275 -765 -241 -731
rect -275 -833 -241 -799
rect -275 -901 -241 -867
rect -275 -969 -241 -935
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect 241 935 275 969
rect 241 867 275 901
rect 241 799 275 833
rect 241 731 275 765
rect 241 663 275 697
rect 241 595 275 629
rect 241 527 275 561
rect 241 459 275 493
rect 241 391 275 425
rect 241 323 275 357
rect 241 255 275 289
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect 241 -289 275 -255
rect 241 -357 275 -323
rect 241 -425 275 -391
rect 241 -493 275 -459
rect 241 -561 275 -527
rect 241 -629 275 -595
rect 241 -697 275 -663
rect 241 -765 275 -731
rect 241 -833 275 -799
rect 241 -901 275 -867
rect 241 -969 275 -935
rect 499 935 533 969
rect 499 867 533 901
rect 499 799 533 833
rect 499 731 533 765
rect 499 663 533 697
rect 499 595 533 629
rect 499 527 533 561
rect 499 459 533 493
rect 499 391 533 425
rect 499 323 533 357
rect 499 255 533 289
rect 499 187 533 221
rect 499 119 533 153
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 499 -153 533 -119
rect 499 -221 533 -187
rect 499 -289 533 -255
rect 499 -357 533 -323
rect 499 -425 533 -391
rect 499 -493 533 -459
rect 499 -561 533 -527
rect 499 -629 533 -595
rect 499 -697 533 -663
rect 499 -765 533 -731
rect 499 -833 533 -799
rect 499 -901 533 -867
rect 499 -969 533 -935
<< psubdiff >>
rect -647 1140 -527 1174
rect -493 1140 -459 1174
rect -425 1140 -391 1174
rect -357 1140 -323 1174
rect -289 1140 -255 1174
rect -221 1140 -187 1174
rect -153 1140 -119 1174
rect -85 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 85 1174
rect 119 1140 153 1174
rect 187 1140 221 1174
rect 255 1140 289 1174
rect 323 1140 357 1174
rect 391 1140 425 1174
rect 459 1140 493 1174
rect 527 1140 647 1174
rect -647 1071 -613 1140
rect -647 1003 -613 1037
rect 613 1071 647 1140
rect 613 1003 647 1037
rect -647 935 -613 969
rect -647 867 -613 901
rect -647 799 -613 833
rect -647 731 -613 765
rect -647 663 -613 697
rect -647 595 -613 629
rect -647 527 -613 561
rect -647 459 -613 493
rect -647 391 -613 425
rect -647 323 -613 357
rect -647 255 -613 289
rect -647 187 -613 221
rect -647 119 -613 153
rect -647 51 -613 85
rect -647 -17 -613 17
rect -647 -85 -613 -51
rect -647 -153 -613 -119
rect -647 -221 -613 -187
rect -647 -289 -613 -255
rect -647 -357 -613 -323
rect -647 -425 -613 -391
rect -647 -493 -613 -459
rect -647 -561 -613 -527
rect -647 -629 -613 -595
rect -647 -697 -613 -663
rect -647 -765 -613 -731
rect -647 -833 -613 -799
rect -647 -901 -613 -867
rect -647 -969 -613 -935
rect 613 935 647 969
rect 613 867 647 901
rect 613 799 647 833
rect 613 731 647 765
rect 613 663 647 697
rect 613 595 647 629
rect 613 527 647 561
rect 613 459 647 493
rect 613 391 647 425
rect 613 323 647 357
rect 613 255 647 289
rect 613 187 647 221
rect 613 119 647 153
rect 613 51 647 85
rect 613 -17 647 17
rect 613 -85 647 -51
rect 613 -153 647 -119
rect 613 -221 647 -187
rect 613 -289 647 -255
rect 613 -357 647 -323
rect 613 -425 647 -391
rect 613 -493 647 -459
rect 613 -561 647 -527
rect 613 -629 647 -595
rect 613 -697 647 -663
rect 613 -765 647 -731
rect 613 -833 647 -799
rect 613 -901 647 -867
rect 613 -969 647 -935
rect -647 -1037 -613 -1003
rect -647 -1140 -613 -1071
rect 613 -1037 647 -1003
rect 613 -1140 647 -1071
rect -647 -1174 -527 -1140
rect -493 -1174 -459 -1140
rect -425 -1174 -391 -1140
rect -357 -1174 -323 -1140
rect -289 -1174 -255 -1140
rect -221 -1174 -187 -1140
rect -153 -1174 -119 -1140
rect -85 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 85 -1140
rect 119 -1174 153 -1140
rect 187 -1174 221 -1140
rect 255 -1174 289 -1140
rect 323 -1174 357 -1140
rect 391 -1174 425 -1140
rect 459 -1174 493 -1140
rect 527 -1174 647 -1140
<< psubdiffcont >>
rect -527 1140 -493 1174
rect -459 1140 -425 1174
rect -391 1140 -357 1174
rect -323 1140 -289 1174
rect -255 1140 -221 1174
rect -187 1140 -153 1174
rect -119 1140 -85 1174
rect -51 1140 -17 1174
rect 17 1140 51 1174
rect 85 1140 119 1174
rect 153 1140 187 1174
rect 221 1140 255 1174
rect 289 1140 323 1174
rect 357 1140 391 1174
rect 425 1140 459 1174
rect 493 1140 527 1174
rect -647 1037 -613 1071
rect -647 969 -613 1003
rect 613 1037 647 1071
rect -647 901 -613 935
rect -647 833 -613 867
rect -647 765 -613 799
rect -647 697 -613 731
rect -647 629 -613 663
rect -647 561 -613 595
rect -647 493 -613 527
rect -647 425 -613 459
rect -647 357 -613 391
rect -647 289 -613 323
rect -647 221 -613 255
rect -647 153 -613 187
rect -647 85 -613 119
rect -647 17 -613 51
rect -647 -51 -613 -17
rect -647 -119 -613 -85
rect -647 -187 -613 -153
rect -647 -255 -613 -221
rect -647 -323 -613 -289
rect -647 -391 -613 -357
rect -647 -459 -613 -425
rect -647 -527 -613 -493
rect -647 -595 -613 -561
rect -647 -663 -613 -629
rect -647 -731 -613 -697
rect -647 -799 -613 -765
rect -647 -867 -613 -833
rect -647 -935 -613 -901
rect -647 -1003 -613 -969
rect 613 969 647 1003
rect 613 901 647 935
rect 613 833 647 867
rect 613 765 647 799
rect 613 697 647 731
rect 613 629 647 663
rect 613 561 647 595
rect 613 493 647 527
rect 613 425 647 459
rect 613 357 647 391
rect 613 289 647 323
rect 613 221 647 255
rect 613 153 647 187
rect 613 85 647 119
rect 613 17 647 51
rect 613 -51 647 -17
rect 613 -119 647 -85
rect 613 -187 647 -153
rect 613 -255 647 -221
rect 613 -323 647 -289
rect 613 -391 647 -357
rect 613 -459 647 -425
rect 613 -527 647 -493
rect 613 -595 647 -561
rect 613 -663 647 -629
rect 613 -731 647 -697
rect 613 -799 647 -765
rect 613 -867 647 -833
rect 613 -935 647 -901
rect -647 -1071 -613 -1037
rect 613 -1003 647 -969
rect 613 -1071 647 -1037
rect -527 -1174 -493 -1140
rect -459 -1174 -425 -1140
rect -391 -1174 -357 -1140
rect -323 -1174 -289 -1140
rect -255 -1174 -221 -1140
rect -187 -1174 -153 -1140
rect -119 -1174 -85 -1140
rect -51 -1174 -17 -1140
rect 17 -1174 51 -1140
rect 85 -1174 119 -1140
rect 153 -1174 187 -1140
rect 221 -1174 255 -1140
rect 289 -1174 323 -1140
rect 357 -1174 391 -1140
rect 425 -1174 459 -1140
rect 493 -1174 527 -1140
<< poly >>
rect -487 1072 -287 1088
rect -487 1038 -438 1072
rect -404 1038 -370 1072
rect -336 1038 -287 1072
rect -487 1000 -287 1038
rect -229 1072 -29 1088
rect -229 1038 -180 1072
rect -146 1038 -112 1072
rect -78 1038 -29 1072
rect -229 1000 -29 1038
rect 29 1072 229 1088
rect 29 1038 78 1072
rect 112 1038 146 1072
rect 180 1038 229 1072
rect 29 1000 229 1038
rect 287 1072 487 1088
rect 287 1038 336 1072
rect 370 1038 404 1072
rect 438 1038 487 1072
rect 287 1000 487 1038
rect -487 -1038 -287 -1000
rect -487 -1072 -438 -1038
rect -404 -1072 -370 -1038
rect -336 -1072 -287 -1038
rect -487 -1088 -287 -1072
rect -229 -1038 -29 -1000
rect -229 -1072 -180 -1038
rect -146 -1072 -112 -1038
rect -78 -1072 -29 -1038
rect -229 -1088 -29 -1072
rect 29 -1038 229 -1000
rect 29 -1072 78 -1038
rect 112 -1072 146 -1038
rect 180 -1072 229 -1038
rect 29 -1088 229 -1072
rect 287 -1038 487 -1000
rect 287 -1072 336 -1038
rect 370 -1072 404 -1038
rect 438 -1072 487 -1038
rect 287 -1088 487 -1072
<< polycont >>
rect -438 1038 -404 1072
rect -370 1038 -336 1072
rect -180 1038 -146 1072
rect -112 1038 -78 1072
rect 78 1038 112 1072
rect 146 1038 180 1072
rect 336 1038 370 1072
rect 404 1038 438 1072
rect -438 -1072 -404 -1038
rect -370 -1072 -336 -1038
rect -180 -1072 -146 -1038
rect -112 -1072 -78 -1038
rect 78 -1072 112 -1038
rect 146 -1072 180 -1038
rect 336 -1072 370 -1038
rect 404 -1072 438 -1038
<< locali >>
rect -647 1140 -527 1174
rect -493 1140 -459 1174
rect -425 1140 -391 1174
rect -357 1140 -323 1174
rect -289 1140 -255 1174
rect -221 1140 -187 1174
rect -153 1140 -119 1174
rect -85 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 85 1174
rect 119 1140 153 1174
rect 187 1140 221 1174
rect 255 1140 289 1174
rect 323 1140 357 1174
rect 391 1140 425 1174
rect 459 1140 493 1174
rect 527 1140 647 1174
rect -647 1071 -613 1140
rect -487 1038 -440 1072
rect -404 1038 -370 1072
rect -334 1038 -287 1072
rect -229 1038 -182 1072
rect -146 1038 -112 1072
rect -76 1038 -29 1072
rect 29 1038 76 1072
rect 112 1038 146 1072
rect 182 1038 229 1072
rect 287 1038 334 1072
rect 370 1038 404 1072
rect 440 1038 487 1072
rect 613 1071 647 1140
rect -647 1003 -613 1037
rect -647 935 -613 969
rect -647 867 -613 901
rect -647 799 -613 833
rect -647 731 -613 765
rect -647 663 -613 697
rect -647 595 -613 629
rect -647 527 -613 561
rect -647 459 -613 493
rect -647 391 -613 425
rect -647 323 -613 357
rect -647 255 -613 289
rect -647 187 -613 221
rect -647 119 -613 153
rect -647 51 -613 85
rect -647 -17 -613 17
rect -647 -85 -613 -51
rect -647 -153 -613 -119
rect -647 -221 -613 -187
rect -647 -289 -613 -255
rect -647 -357 -613 -323
rect -647 -425 -613 -391
rect -647 -493 -613 -459
rect -647 -561 -613 -527
rect -647 -629 -613 -595
rect -647 -697 -613 -663
rect -647 -765 -613 -731
rect -647 -833 -613 -799
rect -647 -901 -613 -867
rect -647 -969 -613 -935
rect -647 -1037 -613 -1003
rect -533 969 -499 1004
rect -533 901 -499 919
rect -533 833 -499 847
rect -533 765 -499 775
rect -533 697 -499 703
rect -533 629 -499 631
rect -533 593 -499 595
rect -533 521 -499 527
rect -533 449 -499 459
rect -533 377 -499 391
rect -533 305 -499 323
rect -533 233 -499 255
rect -533 161 -499 187
rect -533 89 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -89
rect -533 -187 -499 -161
rect -533 -255 -499 -233
rect -533 -323 -499 -305
rect -533 -391 -499 -377
rect -533 -459 -499 -449
rect -533 -527 -499 -521
rect -533 -595 -499 -593
rect -533 -631 -499 -629
rect -533 -703 -499 -697
rect -533 -775 -499 -765
rect -533 -847 -499 -833
rect -533 -919 -499 -901
rect -533 -1004 -499 -969
rect -275 969 -241 1004
rect -275 901 -241 919
rect -275 833 -241 847
rect -275 765 -241 775
rect -275 697 -241 703
rect -275 629 -241 631
rect -275 593 -241 595
rect -275 521 -241 527
rect -275 449 -241 459
rect -275 377 -241 391
rect -275 305 -241 323
rect -275 233 -241 255
rect -275 161 -241 187
rect -275 89 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -89
rect -275 -187 -241 -161
rect -275 -255 -241 -233
rect -275 -323 -241 -305
rect -275 -391 -241 -377
rect -275 -459 -241 -449
rect -275 -527 -241 -521
rect -275 -595 -241 -593
rect -275 -631 -241 -629
rect -275 -703 -241 -697
rect -275 -775 -241 -765
rect -275 -847 -241 -833
rect -275 -919 -241 -901
rect -275 -1004 -241 -969
rect -17 969 17 1004
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -1004 17 -969
rect 241 969 275 1004
rect 241 901 275 919
rect 241 833 275 847
rect 241 765 275 775
rect 241 697 275 703
rect 241 629 275 631
rect 241 593 275 595
rect 241 521 275 527
rect 241 449 275 459
rect 241 377 275 391
rect 241 305 275 323
rect 241 233 275 255
rect 241 161 275 187
rect 241 89 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -89
rect 241 -187 275 -161
rect 241 -255 275 -233
rect 241 -323 275 -305
rect 241 -391 275 -377
rect 241 -459 275 -449
rect 241 -527 275 -521
rect 241 -595 275 -593
rect 241 -631 275 -629
rect 241 -703 275 -697
rect 241 -775 275 -765
rect 241 -847 275 -833
rect 241 -919 275 -901
rect 241 -1004 275 -969
rect 499 969 533 1004
rect 499 901 533 919
rect 499 833 533 847
rect 499 765 533 775
rect 499 697 533 703
rect 499 629 533 631
rect 499 593 533 595
rect 499 521 533 527
rect 499 449 533 459
rect 499 377 533 391
rect 499 305 533 323
rect 499 233 533 255
rect 499 161 533 187
rect 499 89 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -89
rect 499 -187 533 -161
rect 499 -255 533 -233
rect 499 -323 533 -305
rect 499 -391 533 -377
rect 499 -459 533 -449
rect 499 -527 533 -521
rect 499 -595 533 -593
rect 499 -631 533 -629
rect 499 -703 533 -697
rect 499 -775 533 -765
rect 499 -847 533 -833
rect 499 -919 533 -901
rect 499 -1004 533 -969
rect 613 1003 647 1037
rect 613 935 647 969
rect 613 867 647 901
rect 613 799 647 833
rect 613 731 647 765
rect 613 663 647 697
rect 613 595 647 629
rect 613 527 647 561
rect 613 459 647 493
rect 613 391 647 425
rect 613 323 647 357
rect 613 255 647 289
rect 613 187 647 221
rect 613 119 647 153
rect 613 51 647 85
rect 613 -17 647 17
rect 613 -85 647 -51
rect 613 -153 647 -119
rect 613 -221 647 -187
rect 613 -289 647 -255
rect 613 -357 647 -323
rect 613 -425 647 -391
rect 613 -493 647 -459
rect 613 -561 647 -527
rect 613 -629 647 -595
rect 613 -697 647 -663
rect 613 -765 647 -731
rect 613 -833 647 -799
rect 613 -901 647 -867
rect 613 -969 647 -935
rect 613 -1037 647 -1003
rect -647 -1140 -613 -1071
rect -487 -1072 -440 -1038
rect -404 -1072 -370 -1038
rect -334 -1072 -287 -1038
rect -229 -1072 -182 -1038
rect -146 -1072 -112 -1038
rect -76 -1072 -29 -1038
rect 29 -1072 76 -1038
rect 112 -1072 146 -1038
rect 182 -1072 229 -1038
rect 287 -1072 334 -1038
rect 370 -1072 404 -1038
rect 440 -1072 487 -1038
rect 613 -1140 647 -1071
rect -647 -1174 -527 -1140
rect -493 -1174 -459 -1140
rect -425 -1174 -391 -1140
rect -357 -1174 -323 -1140
rect -289 -1174 -255 -1140
rect -221 -1174 -187 -1140
rect -153 -1174 -119 -1140
rect -85 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 85 -1140
rect 119 -1174 153 -1140
rect 187 -1174 221 -1140
rect 255 -1174 289 -1140
rect 323 -1174 357 -1140
rect 391 -1174 425 -1140
rect 459 -1174 493 -1140
rect 527 -1174 647 -1140
<< viali >>
rect -440 1038 -438 1072
rect -438 1038 -406 1072
rect -368 1038 -336 1072
rect -336 1038 -334 1072
rect -182 1038 -180 1072
rect -180 1038 -148 1072
rect -110 1038 -78 1072
rect -78 1038 -76 1072
rect 76 1038 78 1072
rect 78 1038 110 1072
rect 148 1038 180 1072
rect 180 1038 182 1072
rect 334 1038 336 1072
rect 336 1038 368 1072
rect 406 1038 438 1072
rect 438 1038 440 1072
rect -533 935 -499 953
rect -533 919 -499 935
rect -533 867 -499 881
rect -533 847 -499 867
rect -533 799 -499 809
rect -533 775 -499 799
rect -533 731 -499 737
rect -533 703 -499 731
rect -533 663 -499 665
rect -533 631 -499 663
rect -533 561 -499 593
rect -533 559 -499 561
rect -533 493 -499 521
rect -533 487 -499 493
rect -533 425 -499 449
rect -533 415 -499 425
rect -533 357 -499 377
rect -533 343 -499 357
rect -533 289 -499 305
rect -533 271 -499 289
rect -533 221 -499 233
rect -533 199 -499 221
rect -533 153 -499 161
rect -533 127 -499 153
rect -533 85 -499 89
rect -533 55 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -55
rect -533 -89 -499 -85
rect -533 -153 -499 -127
rect -533 -161 -499 -153
rect -533 -221 -499 -199
rect -533 -233 -499 -221
rect -533 -289 -499 -271
rect -533 -305 -499 -289
rect -533 -357 -499 -343
rect -533 -377 -499 -357
rect -533 -425 -499 -415
rect -533 -449 -499 -425
rect -533 -493 -499 -487
rect -533 -521 -499 -493
rect -533 -561 -499 -559
rect -533 -593 -499 -561
rect -533 -663 -499 -631
rect -533 -665 -499 -663
rect -533 -731 -499 -703
rect -533 -737 -499 -731
rect -533 -799 -499 -775
rect -533 -809 -499 -799
rect -533 -867 -499 -847
rect -533 -881 -499 -867
rect -533 -935 -499 -919
rect -533 -953 -499 -935
rect -275 935 -241 953
rect -275 919 -241 935
rect -275 867 -241 881
rect -275 847 -241 867
rect -275 799 -241 809
rect -275 775 -241 799
rect -275 731 -241 737
rect -275 703 -241 731
rect -275 663 -241 665
rect -275 631 -241 663
rect -275 561 -241 593
rect -275 559 -241 561
rect -275 493 -241 521
rect -275 487 -241 493
rect -275 425 -241 449
rect -275 415 -241 425
rect -275 357 -241 377
rect -275 343 -241 357
rect -275 289 -241 305
rect -275 271 -241 289
rect -275 221 -241 233
rect -275 199 -241 221
rect -275 153 -241 161
rect -275 127 -241 153
rect -275 85 -241 89
rect -275 55 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -55
rect -275 -89 -241 -85
rect -275 -153 -241 -127
rect -275 -161 -241 -153
rect -275 -221 -241 -199
rect -275 -233 -241 -221
rect -275 -289 -241 -271
rect -275 -305 -241 -289
rect -275 -357 -241 -343
rect -275 -377 -241 -357
rect -275 -425 -241 -415
rect -275 -449 -241 -425
rect -275 -493 -241 -487
rect -275 -521 -241 -493
rect -275 -561 -241 -559
rect -275 -593 -241 -561
rect -275 -663 -241 -631
rect -275 -665 -241 -663
rect -275 -731 -241 -703
rect -275 -737 -241 -731
rect -275 -799 -241 -775
rect -275 -809 -241 -799
rect -275 -867 -241 -847
rect -275 -881 -241 -867
rect -275 -935 -241 -919
rect -275 -953 -241 -935
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect 241 935 275 953
rect 241 919 275 935
rect 241 867 275 881
rect 241 847 275 867
rect 241 799 275 809
rect 241 775 275 799
rect 241 731 275 737
rect 241 703 275 731
rect 241 663 275 665
rect 241 631 275 663
rect 241 561 275 593
rect 241 559 275 561
rect 241 493 275 521
rect 241 487 275 493
rect 241 425 275 449
rect 241 415 275 425
rect 241 357 275 377
rect 241 343 275 357
rect 241 289 275 305
rect 241 271 275 289
rect 241 221 275 233
rect 241 199 275 221
rect 241 153 275 161
rect 241 127 275 153
rect 241 85 275 89
rect 241 55 275 85
rect 241 -17 275 17
rect 241 -85 275 -55
rect 241 -89 275 -85
rect 241 -153 275 -127
rect 241 -161 275 -153
rect 241 -221 275 -199
rect 241 -233 275 -221
rect 241 -289 275 -271
rect 241 -305 275 -289
rect 241 -357 275 -343
rect 241 -377 275 -357
rect 241 -425 275 -415
rect 241 -449 275 -425
rect 241 -493 275 -487
rect 241 -521 275 -493
rect 241 -561 275 -559
rect 241 -593 275 -561
rect 241 -663 275 -631
rect 241 -665 275 -663
rect 241 -731 275 -703
rect 241 -737 275 -731
rect 241 -799 275 -775
rect 241 -809 275 -799
rect 241 -867 275 -847
rect 241 -881 275 -867
rect 241 -935 275 -919
rect 241 -953 275 -935
rect 499 935 533 953
rect 499 919 533 935
rect 499 867 533 881
rect 499 847 533 867
rect 499 799 533 809
rect 499 775 533 799
rect 499 731 533 737
rect 499 703 533 731
rect 499 663 533 665
rect 499 631 533 663
rect 499 561 533 593
rect 499 559 533 561
rect 499 493 533 521
rect 499 487 533 493
rect 499 425 533 449
rect 499 415 533 425
rect 499 357 533 377
rect 499 343 533 357
rect 499 289 533 305
rect 499 271 533 289
rect 499 221 533 233
rect 499 199 533 221
rect 499 153 533 161
rect 499 127 533 153
rect 499 85 533 89
rect 499 55 533 85
rect 499 -17 533 17
rect 499 -85 533 -55
rect 499 -89 533 -85
rect 499 -153 533 -127
rect 499 -161 533 -153
rect 499 -221 533 -199
rect 499 -233 533 -221
rect 499 -289 533 -271
rect 499 -305 533 -289
rect 499 -357 533 -343
rect 499 -377 533 -357
rect 499 -425 533 -415
rect 499 -449 533 -425
rect 499 -493 533 -487
rect 499 -521 533 -493
rect 499 -561 533 -559
rect 499 -593 533 -561
rect 499 -663 533 -631
rect 499 -665 533 -663
rect 499 -731 533 -703
rect 499 -737 533 -731
rect 499 -799 533 -775
rect 499 -809 533 -799
rect 499 -867 533 -847
rect 499 -881 533 -867
rect 499 -935 533 -919
rect 499 -953 533 -935
rect -440 -1072 -438 -1038
rect -438 -1072 -406 -1038
rect -368 -1072 -336 -1038
rect -336 -1072 -334 -1038
rect -182 -1072 -180 -1038
rect -180 -1072 -148 -1038
rect -110 -1072 -78 -1038
rect -78 -1072 -76 -1038
rect 76 -1072 78 -1038
rect 78 -1072 110 -1038
rect 148 -1072 180 -1038
rect 180 -1072 182 -1038
rect 334 -1072 336 -1038
rect 336 -1072 368 -1038
rect 406 -1072 438 -1038
rect 438 -1072 440 -1038
<< metal1 >>
rect -483 1072 -291 1078
rect -483 1038 -440 1072
rect -406 1038 -368 1072
rect -334 1038 -291 1072
rect -483 1032 -291 1038
rect -225 1072 -33 1078
rect -225 1038 -182 1072
rect -148 1038 -110 1072
rect -76 1038 -33 1072
rect -225 1032 -33 1038
rect 33 1072 225 1078
rect 33 1038 76 1072
rect 110 1038 148 1072
rect 182 1038 225 1072
rect 33 1032 225 1038
rect 291 1072 483 1078
rect 291 1038 334 1072
rect 368 1038 406 1072
rect 440 1038 483 1072
rect 291 1032 483 1038
rect -539 953 -493 1000
rect -539 919 -533 953
rect -499 919 -493 953
rect -539 881 -493 919
rect -539 847 -533 881
rect -499 847 -493 881
rect -539 809 -493 847
rect -539 775 -533 809
rect -499 775 -493 809
rect -539 737 -493 775
rect -539 703 -533 737
rect -499 703 -493 737
rect -539 665 -493 703
rect -539 631 -533 665
rect -499 631 -493 665
rect -539 593 -493 631
rect -539 559 -533 593
rect -499 559 -493 593
rect -539 521 -493 559
rect -539 487 -533 521
rect -499 487 -493 521
rect -539 449 -493 487
rect -539 415 -533 449
rect -499 415 -493 449
rect -539 377 -493 415
rect -539 343 -533 377
rect -499 343 -493 377
rect -539 305 -493 343
rect -539 271 -533 305
rect -499 271 -493 305
rect -539 233 -493 271
rect -539 199 -533 233
rect -499 199 -493 233
rect -539 161 -493 199
rect -539 127 -533 161
rect -499 127 -493 161
rect -539 89 -493 127
rect -539 55 -533 89
rect -499 55 -493 89
rect -539 17 -493 55
rect -539 -17 -533 17
rect -499 -17 -493 17
rect -539 -55 -493 -17
rect -539 -89 -533 -55
rect -499 -89 -493 -55
rect -539 -127 -493 -89
rect -539 -161 -533 -127
rect -499 -161 -493 -127
rect -539 -199 -493 -161
rect -539 -233 -533 -199
rect -499 -233 -493 -199
rect -539 -271 -493 -233
rect -539 -305 -533 -271
rect -499 -305 -493 -271
rect -539 -343 -493 -305
rect -539 -377 -533 -343
rect -499 -377 -493 -343
rect -539 -415 -493 -377
rect -539 -449 -533 -415
rect -499 -449 -493 -415
rect -539 -487 -493 -449
rect -539 -521 -533 -487
rect -499 -521 -493 -487
rect -539 -559 -493 -521
rect -539 -593 -533 -559
rect -499 -593 -493 -559
rect -539 -631 -493 -593
rect -539 -665 -533 -631
rect -499 -665 -493 -631
rect -539 -703 -493 -665
rect -539 -737 -533 -703
rect -499 -737 -493 -703
rect -539 -775 -493 -737
rect -539 -809 -533 -775
rect -499 -809 -493 -775
rect -539 -847 -493 -809
rect -539 -881 -533 -847
rect -499 -881 -493 -847
rect -539 -919 -493 -881
rect -539 -953 -533 -919
rect -499 -953 -493 -919
rect -539 -1000 -493 -953
rect -281 953 -235 1000
rect -281 919 -275 953
rect -241 919 -235 953
rect -281 881 -235 919
rect -281 847 -275 881
rect -241 847 -235 881
rect -281 809 -235 847
rect -281 775 -275 809
rect -241 775 -235 809
rect -281 737 -235 775
rect -281 703 -275 737
rect -241 703 -235 737
rect -281 665 -235 703
rect -281 631 -275 665
rect -241 631 -235 665
rect -281 593 -235 631
rect -281 559 -275 593
rect -241 559 -235 593
rect -281 521 -235 559
rect -281 487 -275 521
rect -241 487 -235 521
rect -281 449 -235 487
rect -281 415 -275 449
rect -241 415 -235 449
rect -281 377 -235 415
rect -281 343 -275 377
rect -241 343 -235 377
rect -281 305 -235 343
rect -281 271 -275 305
rect -241 271 -235 305
rect -281 233 -235 271
rect -281 199 -275 233
rect -241 199 -235 233
rect -281 161 -235 199
rect -281 127 -275 161
rect -241 127 -235 161
rect -281 89 -235 127
rect -281 55 -275 89
rect -241 55 -235 89
rect -281 17 -235 55
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -127 -235 -89
rect -281 -161 -275 -127
rect -241 -161 -235 -127
rect -281 -199 -235 -161
rect -281 -233 -275 -199
rect -241 -233 -235 -199
rect -281 -271 -235 -233
rect -281 -305 -275 -271
rect -241 -305 -235 -271
rect -281 -343 -235 -305
rect -281 -377 -275 -343
rect -241 -377 -235 -343
rect -281 -415 -235 -377
rect -281 -449 -275 -415
rect -241 -449 -235 -415
rect -281 -487 -235 -449
rect -281 -521 -275 -487
rect -241 -521 -235 -487
rect -281 -559 -235 -521
rect -281 -593 -275 -559
rect -241 -593 -235 -559
rect -281 -631 -235 -593
rect -281 -665 -275 -631
rect -241 -665 -235 -631
rect -281 -703 -235 -665
rect -281 -737 -275 -703
rect -241 -737 -235 -703
rect -281 -775 -235 -737
rect -281 -809 -275 -775
rect -241 -809 -235 -775
rect -281 -847 -235 -809
rect -281 -881 -275 -847
rect -241 -881 -235 -847
rect -281 -919 -235 -881
rect -281 -953 -275 -919
rect -241 -953 -235 -919
rect -281 -1000 -235 -953
rect -23 953 23 1000
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -1000 23 -953
rect 235 953 281 1000
rect 235 919 241 953
rect 275 919 281 953
rect 235 881 281 919
rect 235 847 241 881
rect 275 847 281 881
rect 235 809 281 847
rect 235 775 241 809
rect 275 775 281 809
rect 235 737 281 775
rect 235 703 241 737
rect 275 703 281 737
rect 235 665 281 703
rect 235 631 241 665
rect 275 631 281 665
rect 235 593 281 631
rect 235 559 241 593
rect 275 559 281 593
rect 235 521 281 559
rect 235 487 241 521
rect 275 487 281 521
rect 235 449 281 487
rect 235 415 241 449
rect 275 415 281 449
rect 235 377 281 415
rect 235 343 241 377
rect 275 343 281 377
rect 235 305 281 343
rect 235 271 241 305
rect 275 271 281 305
rect 235 233 281 271
rect 235 199 241 233
rect 275 199 281 233
rect 235 161 281 199
rect 235 127 241 161
rect 275 127 281 161
rect 235 89 281 127
rect 235 55 241 89
rect 275 55 281 89
rect 235 17 281 55
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -127 281 -89
rect 235 -161 241 -127
rect 275 -161 281 -127
rect 235 -199 281 -161
rect 235 -233 241 -199
rect 275 -233 281 -199
rect 235 -271 281 -233
rect 235 -305 241 -271
rect 275 -305 281 -271
rect 235 -343 281 -305
rect 235 -377 241 -343
rect 275 -377 281 -343
rect 235 -415 281 -377
rect 235 -449 241 -415
rect 275 -449 281 -415
rect 235 -487 281 -449
rect 235 -521 241 -487
rect 275 -521 281 -487
rect 235 -559 281 -521
rect 235 -593 241 -559
rect 275 -593 281 -559
rect 235 -631 281 -593
rect 235 -665 241 -631
rect 275 -665 281 -631
rect 235 -703 281 -665
rect 235 -737 241 -703
rect 275 -737 281 -703
rect 235 -775 281 -737
rect 235 -809 241 -775
rect 275 -809 281 -775
rect 235 -847 281 -809
rect 235 -881 241 -847
rect 275 -881 281 -847
rect 235 -919 281 -881
rect 235 -953 241 -919
rect 275 -953 281 -919
rect 235 -1000 281 -953
rect 493 953 539 1000
rect 493 919 499 953
rect 533 919 539 953
rect 493 881 539 919
rect 493 847 499 881
rect 533 847 539 881
rect 493 809 539 847
rect 493 775 499 809
rect 533 775 539 809
rect 493 737 539 775
rect 493 703 499 737
rect 533 703 539 737
rect 493 665 539 703
rect 493 631 499 665
rect 533 631 539 665
rect 493 593 539 631
rect 493 559 499 593
rect 533 559 539 593
rect 493 521 539 559
rect 493 487 499 521
rect 533 487 539 521
rect 493 449 539 487
rect 493 415 499 449
rect 533 415 539 449
rect 493 377 539 415
rect 493 343 499 377
rect 533 343 539 377
rect 493 305 539 343
rect 493 271 499 305
rect 533 271 539 305
rect 493 233 539 271
rect 493 199 499 233
rect 533 199 539 233
rect 493 161 539 199
rect 493 127 499 161
rect 533 127 539 161
rect 493 89 539 127
rect 493 55 499 89
rect 533 55 539 89
rect 493 17 539 55
rect 493 -17 499 17
rect 533 -17 539 17
rect 493 -55 539 -17
rect 493 -89 499 -55
rect 533 -89 539 -55
rect 493 -127 539 -89
rect 493 -161 499 -127
rect 533 -161 539 -127
rect 493 -199 539 -161
rect 493 -233 499 -199
rect 533 -233 539 -199
rect 493 -271 539 -233
rect 493 -305 499 -271
rect 533 -305 539 -271
rect 493 -343 539 -305
rect 493 -377 499 -343
rect 533 -377 539 -343
rect 493 -415 539 -377
rect 493 -449 499 -415
rect 533 -449 539 -415
rect 493 -487 539 -449
rect 493 -521 499 -487
rect 533 -521 539 -487
rect 493 -559 539 -521
rect 493 -593 499 -559
rect 533 -593 539 -559
rect 493 -631 539 -593
rect 493 -665 499 -631
rect 533 -665 539 -631
rect 493 -703 539 -665
rect 493 -737 499 -703
rect 533 -737 539 -703
rect 493 -775 539 -737
rect 493 -809 499 -775
rect 533 -809 539 -775
rect 493 -847 539 -809
rect 493 -881 499 -847
rect 533 -881 539 -847
rect 493 -919 539 -881
rect 493 -953 499 -919
rect 533 -953 539 -919
rect 493 -1000 539 -953
rect -483 -1038 -291 -1032
rect -483 -1072 -440 -1038
rect -406 -1072 -368 -1038
rect -334 -1072 -291 -1038
rect -483 -1078 -291 -1072
rect -225 -1038 -33 -1032
rect -225 -1072 -182 -1038
rect -148 -1072 -110 -1038
rect -76 -1072 -33 -1038
rect -225 -1078 -33 -1072
rect 33 -1038 225 -1032
rect 33 -1072 76 -1038
rect 110 -1072 148 -1038
rect 182 -1072 225 -1038
rect 33 -1078 225 -1072
rect 291 -1038 483 -1032
rect 291 -1072 334 -1038
rect 368 -1072 406 -1038
rect 440 -1072 483 -1038
rect 291 -1078 483 -1072
<< properties >>
string FIXED_BBOX -630 -1157 630 1157
<< end >>
