magic
tech sky130A
magscale 1 1
timestamp 1737500400
<< checkpaint >>
rect 0 0 2236 1720
<< locali >>
rect 8 8 2228 64
rect 64 8 2172 64
rect 8 8 2228 64
rect 64 1656 2172 1712
rect 8 1656 2228 1712
rect 8 64 64 1656
rect 8 8 64 1712
rect 2172 64 2228 1656
rect 2172 8 2228 1712
rect 8 8 2228 64
rect 1910 1460 2054 1580
rect 182 1460 326 1580
<< ptapc >>
rect 78 16 118 56
rect 118 16 158 56
rect 158 16 198 56
rect 198 16 238 56
rect 238 16 278 56
rect 278 16 318 56
rect 318 16 358 56
rect 358 16 398 56
rect 398 16 438 56
rect 438 16 478 56
rect 478 16 518 56
rect 518 16 558 56
rect 558 16 598 56
rect 598 16 638 56
rect 638 16 678 56
rect 678 16 718 56
rect 718 16 758 56
rect 758 16 798 56
rect 798 16 838 56
rect 838 16 878 56
rect 878 16 918 56
rect 918 16 958 56
rect 958 16 998 56
rect 998 16 1038 56
rect 1038 16 1078 56
rect 1078 16 1118 56
rect 1118 16 1158 56
rect 1158 16 1198 56
rect 1198 16 1238 56
rect 1238 16 1278 56
rect 1278 16 1318 56
rect 1318 16 1358 56
rect 1358 16 1398 56
rect 1398 16 1438 56
rect 1438 16 1478 56
rect 1478 16 1518 56
rect 1518 16 1558 56
rect 1558 16 1598 56
rect 1598 16 1638 56
rect 1638 16 1678 56
rect 1678 16 1718 56
rect 1718 16 1758 56
rect 1758 16 1798 56
rect 1798 16 1838 56
rect 1838 16 1878 56
rect 1878 16 1918 56
rect 1918 16 1958 56
rect 1958 16 1998 56
rect 1998 16 2038 56
rect 2038 16 2078 56
rect 2078 16 2118 56
rect 2118 16 2158 56
rect 78 1664 118 1704
rect 118 1664 158 1704
rect 158 1664 198 1704
rect 198 1664 238 1704
rect 238 1664 278 1704
rect 278 1664 318 1704
rect 318 1664 358 1704
rect 358 1664 398 1704
rect 398 1664 438 1704
rect 438 1664 478 1704
rect 478 1664 518 1704
rect 518 1664 558 1704
rect 558 1664 598 1704
rect 598 1664 638 1704
rect 638 1664 678 1704
rect 678 1664 718 1704
rect 718 1664 758 1704
rect 758 1664 798 1704
rect 798 1664 838 1704
rect 838 1664 878 1704
rect 878 1664 918 1704
rect 918 1664 958 1704
rect 958 1664 998 1704
rect 998 1664 1038 1704
rect 1038 1664 1078 1704
rect 1078 1664 1118 1704
rect 1118 1664 1158 1704
rect 1158 1664 1198 1704
rect 1198 1664 1238 1704
rect 1238 1664 1278 1704
rect 1278 1664 1318 1704
rect 1318 1664 1358 1704
rect 1358 1664 1398 1704
rect 1398 1664 1438 1704
rect 1438 1664 1478 1704
rect 1478 1664 1518 1704
rect 1518 1664 1558 1704
rect 1558 1664 1598 1704
rect 1598 1664 1638 1704
rect 1638 1664 1678 1704
rect 1678 1664 1718 1704
rect 1718 1664 1758 1704
rect 1758 1664 1798 1704
rect 1798 1664 1838 1704
rect 1838 1664 1878 1704
rect 1878 1664 1918 1704
rect 1918 1664 1958 1704
rect 1958 1664 1998 1704
rect 1998 1664 2038 1704
rect 2038 1664 2078 1704
rect 2078 1664 2118 1704
rect 2118 1664 2158 1704
rect 16 80 56 120
rect 16 120 56 160
rect 16 160 56 200
rect 16 200 56 240
rect 16 240 56 280
rect 16 280 56 320
rect 16 320 56 360
rect 16 360 56 400
rect 16 400 56 440
rect 16 440 56 480
rect 16 480 56 520
rect 16 520 56 560
rect 16 560 56 600
rect 16 600 56 640
rect 16 640 56 680
rect 16 680 56 720
rect 16 720 56 760
rect 16 760 56 800
rect 16 800 56 840
rect 16 840 56 880
rect 16 880 56 920
rect 16 920 56 960
rect 16 960 56 1000
rect 16 1000 56 1040
rect 16 1040 56 1080
rect 16 1080 56 1120
rect 16 1120 56 1160
rect 16 1160 56 1200
rect 16 1200 56 1240
rect 16 1240 56 1280
rect 16 1280 56 1320
rect 16 1320 56 1360
rect 16 1360 56 1400
rect 16 1400 56 1440
rect 16 1440 56 1480
rect 16 1480 56 1520
rect 16 1520 56 1560
rect 16 1560 56 1600
rect 16 1600 56 1640
rect 2180 80 2220 120
rect 2180 120 2220 160
rect 2180 160 2220 200
rect 2180 200 2220 240
rect 2180 240 2220 280
rect 2180 280 2220 320
rect 2180 320 2220 360
rect 2180 360 2220 400
rect 2180 400 2220 440
rect 2180 440 2220 480
rect 2180 480 2220 520
rect 2180 520 2220 560
rect 2180 560 2220 600
rect 2180 600 2220 640
rect 2180 640 2220 680
rect 2180 680 2220 720
rect 2180 720 2220 760
rect 2180 760 2220 800
rect 2180 800 2220 840
rect 2180 840 2220 880
rect 2180 880 2220 920
rect 2180 920 2220 960
rect 2180 960 2220 1000
rect 2180 1000 2220 1040
rect 2180 1040 2220 1080
rect 2180 1080 2220 1120
rect 2180 1120 2220 1160
rect 2180 1160 2220 1200
rect 2180 1200 2220 1240
rect 2180 1240 2220 1280
rect 2180 1280 2220 1320
rect 2180 1320 2220 1360
rect 2180 1360 2220 1400
rect 2180 1400 2220 1440
rect 2180 1440 2220 1480
rect 2180 1480 2220 1520
rect 2180 1520 2220 1560
rect 2180 1560 2220 1600
rect 2180 1600 2220 1640
<< ptap >>
rect 0 0 2236 72
rect 0 1648 2236 1720
rect 0 0 72 1720
rect 2164 0 2236 1720
use JNWTR_RES16 XA1 
transform 1 0 200 0 1 200
box 200 200 2036 1520
<< labels >>
flabel locali s 8 8 2228 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 1910 1460 2054 1580 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 182 1460 326 1580 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2236 1720
<< end >>
