magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 704 400
<< pdiff >>
rect 208 100 496 140
rect 208 140 496 180
rect 208 180 496 220
rect 208 220 496 260
rect 208 260 496 300
<< ntap >>
rect -48 -20 48 20
rect 656 -20 752 20
rect -48 20 48 60
rect 656 20 752 60
rect -48 60 48 100
rect 656 60 752 100
rect -48 100 48 140
rect 656 100 752 140
rect -48 140 48 180
rect 656 140 752 180
rect -48 180 48 220
rect 656 180 752 220
rect -48 220 48 260
rect 656 220 752 260
rect -48 260 48 300
rect 656 260 752 300
rect -48 300 48 340
rect 656 300 752 340
rect -48 340 48 380
rect 656 340 752 380
rect -48 380 48 420
rect 656 380 752 420
<< poly >>
rect 80 -11 624 11
rect 80 69 624 91
rect 80 149 624 171
rect 80 229 624 251
rect 80 309 624 331
rect 80 389 624 411
rect 80 140 112 180
rect 592 140 624 180
rect 80 180 112 220
rect 592 180 624 220
rect 80 220 112 260
rect 592 220 624 260
<< m1 >>
rect 80 180 112 220
rect 144 300 240 340
rect 464 20 560 60
rect 80 20 112 60
rect 144 20 240 60
rect 464 20 560 60
rect 80 60 112 100
rect 144 60 240 100
rect 464 60 560 100
rect 80 100 112 140
rect 144 100 240 140
rect 464 100 560 140
rect 80 140 112 180
rect 144 140 240 180
rect 464 140 560 180
rect 80 180 112 220
rect 144 180 240 220
rect 464 180 560 220
rect 80 220 112 260
rect 144 220 240 260
rect 464 220 560 260
rect 80 260 112 300
rect 144 260 240 300
rect 464 260 560 300
rect 80 300 112 340
rect 144 300 240 340
rect 464 300 560 340
rect 80 340 112 380
rect 144 340 240 380
rect 464 340 560 380
<< pcontact >>
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 597 150 618 160
rect 597 160 618 170
rect 597 170 618 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 597 180 618 190
rect 597 190 618 200
rect 597 200 618 210
rect 597 210 618 220
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 597 220 618 230
rect 597 230 618 240
rect 597 240 618 250
<< locali >>
rect -48 -20 48 20
rect 656 -20 752 20
rect -48 20 48 60
rect 656 20 752 60
rect -48 60 48 100
rect 656 60 752 100
rect -48 100 48 140
rect 144 100 496 140
rect 656 100 752 140
rect -48 140 48 180
rect 80 140 112 180
rect 592 140 624 180
rect 656 140 752 180
rect -48 180 48 220
rect -48 180 48 220
rect 80 180 112 220
rect 208 180 560 220
rect 592 180 624 220
rect 656 180 752 220
rect -48 220 48 260
rect 80 220 112 260
rect 592 220 624 260
rect 656 220 752 260
rect -48 260 48 300
rect 144 260 496 300
rect 656 260 752 300
rect -48 300 48 340
rect 656 300 752 340
rect -48 340 48 380
rect 656 340 752 380
rect -48 380 48 420
rect 656 380 752 420
<< ntapc >>
rect -16 100 16 140
rect 688 100 720 140
rect -16 140 16 180
rect 688 140 720 180
rect -16 180 16 220
rect 688 180 720 220
rect -16 220 16 260
rect 688 220 720 260
rect -16 260 16 300
rect 688 260 720 300
<< pdcontact >>
rect 224 110 240 120
rect 224 120 240 130
rect 240 110 272 120
rect 240 120 272 130
rect 272 110 304 120
rect 272 120 304 130
rect 304 110 336 120
rect 304 120 336 130
rect 336 110 368 120
rect 336 120 368 130
rect 368 110 400 120
rect 368 120 400 130
rect 400 110 432 120
rect 400 120 432 130
rect 432 110 464 120
rect 432 120 464 130
rect 464 110 480 120
rect 464 120 480 130
rect 224 190 240 200
rect 224 200 240 210
rect 240 190 272 200
rect 240 200 272 210
rect 272 190 304 200
rect 272 200 304 210
rect 304 190 336 200
rect 304 200 336 210
rect 336 190 368 200
rect 336 200 368 210
rect 368 190 400 200
rect 368 200 400 210
rect 400 190 432 200
rect 400 200 432 210
rect 432 190 464 200
rect 432 200 464 210
rect 464 190 480 200
rect 464 200 480 210
rect 224 270 240 280
rect 224 280 240 290
rect 240 270 272 280
rect 240 280 272 290
rect 272 270 304 280
rect 272 280 304 290
rect 304 270 336 280
rect 304 280 336 290
rect 336 270 368 280
rect 336 280 368 290
rect 368 270 400 280
rect 368 280 400 290
rect 400 270 432 280
rect 400 280 432 290
rect 432 270 464 280
rect 432 280 464 290
rect 464 270 480 280
rect 464 280 480 290
<< viali >>
rect 160 104 176 108
rect 160 108 176 112
rect 160 112 176 116
rect 160 116 176 120
rect 160 120 176 124
rect 160 124 176 128
rect 160 128 176 132
rect 160 132 176 136
rect 176 104 208 108
rect 176 108 208 112
rect 176 112 208 116
rect 176 116 208 120
rect 176 120 208 124
rect 176 124 208 128
rect 176 128 208 132
rect 176 132 208 136
rect 208 104 224 108
rect 208 108 224 112
rect 208 112 224 116
rect 208 116 224 120
rect 208 120 224 124
rect 208 124 224 128
rect 208 128 224 132
rect 208 132 224 136
rect 85 150 106 160
rect 85 160 106 170
rect 85 170 106 180
rect 85 180 106 190
rect 85 190 106 200
rect 85 200 106 210
rect 85 210 106 220
rect 480 184 496 188
rect 480 188 496 192
rect 480 192 496 196
rect 480 196 496 200
rect 480 200 496 204
rect 480 204 496 208
rect 480 208 496 212
rect 480 212 496 216
rect 496 184 528 188
rect 496 188 528 192
rect 496 192 528 196
rect 496 196 528 200
rect 496 200 528 204
rect 496 204 528 208
rect 496 208 528 212
rect 496 212 528 216
rect 528 184 544 188
rect 528 188 544 192
rect 528 192 544 196
rect 528 196 544 200
rect 528 200 544 204
rect 528 204 544 208
rect 528 208 544 212
rect 528 212 544 216
rect 85 220 106 230
rect 85 230 106 240
rect 85 240 106 250
rect 160 264 176 268
rect 160 268 176 272
rect 160 272 176 276
rect 160 276 176 280
rect 160 280 176 284
rect 160 284 176 288
rect 160 288 176 292
rect 160 292 176 296
rect 176 264 208 268
rect 176 268 208 272
rect 176 272 208 276
rect 176 276 208 280
rect 176 280 208 284
rect 176 284 208 288
rect 176 288 208 292
rect 176 292 208 296
rect 208 264 224 268
rect 208 268 224 272
rect 208 272 224 276
rect 208 276 224 280
rect 208 280 224 284
rect 208 284 224 288
rect 208 288 224 292
rect 208 292 224 296
<< nwell >>
rect -92 -64 796 464
<< labels >>
flabel m1 s 80 180 112 220 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel m1 s 144 300 240 340 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -48 180 48 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel m1 s 464 20 560 60 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 704 400
<< end >>
