magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -2696 -319 2696 319
<< pmos >>
rect -2500 -100 2500 100
<< pdiff >>
rect -2558 85 -2500 100
rect -2558 51 -2546 85
rect -2512 51 -2500 85
rect -2558 17 -2500 51
rect -2558 -17 -2546 17
rect -2512 -17 -2500 17
rect -2558 -51 -2500 -17
rect -2558 -85 -2546 -51
rect -2512 -85 -2500 -51
rect -2558 -100 -2500 -85
rect 2500 85 2558 100
rect 2500 51 2512 85
rect 2546 51 2558 85
rect 2500 17 2558 51
rect 2500 -17 2512 17
rect 2546 -17 2558 17
rect 2500 -51 2558 -17
rect 2500 -85 2512 -51
rect 2546 -85 2558 -51
rect 2500 -100 2558 -85
<< pdiffc >>
rect -2546 51 -2512 85
rect -2546 -17 -2512 17
rect -2546 -85 -2512 -51
rect 2512 51 2546 85
rect 2512 -17 2546 17
rect 2512 -85 2546 -51
<< nsubdiff >>
rect -2660 249 -2533 283
rect -2499 249 -2465 283
rect -2431 249 -2397 283
rect -2363 249 -2329 283
rect -2295 249 -2261 283
rect -2227 249 -2193 283
rect -2159 249 -2125 283
rect -2091 249 -2057 283
rect -2023 249 -1989 283
rect -1955 249 -1921 283
rect -1887 249 -1853 283
rect -1819 249 -1785 283
rect -1751 249 -1717 283
rect -1683 249 -1649 283
rect -1615 249 -1581 283
rect -1547 249 -1513 283
rect -1479 249 -1445 283
rect -1411 249 -1377 283
rect -1343 249 -1309 283
rect -1275 249 -1241 283
rect -1207 249 -1173 283
rect -1139 249 -1105 283
rect -1071 249 -1037 283
rect -1003 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1003 283
rect 1037 249 1071 283
rect 1105 249 1139 283
rect 1173 249 1207 283
rect 1241 249 1275 283
rect 1309 249 1343 283
rect 1377 249 1411 283
rect 1445 249 1479 283
rect 1513 249 1547 283
rect 1581 249 1615 283
rect 1649 249 1683 283
rect 1717 249 1751 283
rect 1785 249 1819 283
rect 1853 249 1887 283
rect 1921 249 1955 283
rect 1989 249 2023 283
rect 2057 249 2091 283
rect 2125 249 2159 283
rect 2193 249 2227 283
rect 2261 249 2295 283
rect 2329 249 2363 283
rect 2397 249 2431 283
rect 2465 249 2499 283
rect 2533 249 2660 283
rect -2660 187 -2626 249
rect -2660 119 -2626 153
rect 2626 187 2660 249
rect 2626 119 2660 153
rect -2660 51 -2626 85
rect -2660 -17 -2626 17
rect -2660 -85 -2626 -51
rect 2626 51 2660 85
rect 2626 -17 2660 17
rect 2626 -85 2660 -51
rect -2660 -153 -2626 -119
rect -2660 -249 -2626 -187
rect 2626 -153 2660 -119
rect 2626 -249 2660 -187
rect -2660 -283 -2533 -249
rect -2499 -283 -2465 -249
rect -2431 -283 -2397 -249
rect -2363 -283 -2329 -249
rect -2295 -283 -2261 -249
rect -2227 -283 -2193 -249
rect -2159 -283 -2125 -249
rect -2091 -283 -2057 -249
rect -2023 -283 -1989 -249
rect -1955 -283 -1921 -249
rect -1887 -283 -1853 -249
rect -1819 -283 -1785 -249
rect -1751 -283 -1717 -249
rect -1683 -283 -1649 -249
rect -1615 -283 -1581 -249
rect -1547 -283 -1513 -249
rect -1479 -283 -1445 -249
rect -1411 -283 -1377 -249
rect -1343 -283 -1309 -249
rect -1275 -283 -1241 -249
rect -1207 -283 -1173 -249
rect -1139 -283 -1105 -249
rect -1071 -283 -1037 -249
rect -1003 -283 -969 -249
rect -935 -283 -901 -249
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
rect 901 -283 935 -249
rect 969 -283 1003 -249
rect 1037 -283 1071 -249
rect 1105 -283 1139 -249
rect 1173 -283 1207 -249
rect 1241 -283 1275 -249
rect 1309 -283 1343 -249
rect 1377 -283 1411 -249
rect 1445 -283 1479 -249
rect 1513 -283 1547 -249
rect 1581 -283 1615 -249
rect 1649 -283 1683 -249
rect 1717 -283 1751 -249
rect 1785 -283 1819 -249
rect 1853 -283 1887 -249
rect 1921 -283 1955 -249
rect 1989 -283 2023 -249
rect 2057 -283 2091 -249
rect 2125 -283 2159 -249
rect 2193 -283 2227 -249
rect 2261 -283 2295 -249
rect 2329 -283 2363 -249
rect 2397 -283 2431 -249
rect 2465 -283 2499 -249
rect 2533 -283 2660 -249
<< nsubdiffcont >>
rect -2533 249 -2499 283
rect -2465 249 -2431 283
rect -2397 249 -2363 283
rect -2329 249 -2295 283
rect -2261 249 -2227 283
rect -2193 249 -2159 283
rect -2125 249 -2091 283
rect -2057 249 -2023 283
rect -1989 249 -1955 283
rect -1921 249 -1887 283
rect -1853 249 -1819 283
rect -1785 249 -1751 283
rect -1717 249 -1683 283
rect -1649 249 -1615 283
rect -1581 249 -1547 283
rect -1513 249 -1479 283
rect -1445 249 -1411 283
rect -1377 249 -1343 283
rect -1309 249 -1275 283
rect -1241 249 -1207 283
rect -1173 249 -1139 283
rect -1105 249 -1071 283
rect -1037 249 -1003 283
rect -969 249 -935 283
rect -901 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 901 283
rect 935 249 969 283
rect 1003 249 1037 283
rect 1071 249 1105 283
rect 1139 249 1173 283
rect 1207 249 1241 283
rect 1275 249 1309 283
rect 1343 249 1377 283
rect 1411 249 1445 283
rect 1479 249 1513 283
rect 1547 249 1581 283
rect 1615 249 1649 283
rect 1683 249 1717 283
rect 1751 249 1785 283
rect 1819 249 1853 283
rect 1887 249 1921 283
rect 1955 249 1989 283
rect 2023 249 2057 283
rect 2091 249 2125 283
rect 2159 249 2193 283
rect 2227 249 2261 283
rect 2295 249 2329 283
rect 2363 249 2397 283
rect 2431 249 2465 283
rect 2499 249 2533 283
rect -2660 153 -2626 187
rect -2660 85 -2626 119
rect 2626 153 2660 187
rect -2660 17 -2626 51
rect -2660 -51 -2626 -17
rect -2660 -119 -2626 -85
rect 2626 85 2660 119
rect 2626 17 2660 51
rect 2626 -51 2660 -17
rect -2660 -187 -2626 -153
rect 2626 -119 2660 -85
rect 2626 -187 2660 -153
rect -2533 -283 -2499 -249
rect -2465 -283 -2431 -249
rect -2397 -283 -2363 -249
rect -2329 -283 -2295 -249
rect -2261 -283 -2227 -249
rect -2193 -283 -2159 -249
rect -2125 -283 -2091 -249
rect -2057 -283 -2023 -249
rect -1989 -283 -1955 -249
rect -1921 -283 -1887 -249
rect -1853 -283 -1819 -249
rect -1785 -283 -1751 -249
rect -1717 -283 -1683 -249
rect -1649 -283 -1615 -249
rect -1581 -283 -1547 -249
rect -1513 -283 -1479 -249
rect -1445 -283 -1411 -249
rect -1377 -283 -1343 -249
rect -1309 -283 -1275 -249
rect -1241 -283 -1207 -249
rect -1173 -283 -1139 -249
rect -1105 -283 -1071 -249
rect -1037 -283 -1003 -249
rect -969 -283 -935 -249
rect -901 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 901 -249
rect 935 -283 969 -249
rect 1003 -283 1037 -249
rect 1071 -283 1105 -249
rect 1139 -283 1173 -249
rect 1207 -283 1241 -249
rect 1275 -283 1309 -249
rect 1343 -283 1377 -249
rect 1411 -283 1445 -249
rect 1479 -283 1513 -249
rect 1547 -283 1581 -249
rect 1615 -283 1649 -249
rect 1683 -283 1717 -249
rect 1751 -283 1785 -249
rect 1819 -283 1853 -249
rect 1887 -283 1921 -249
rect 1955 -283 1989 -249
rect 2023 -283 2057 -249
rect 2091 -283 2125 -249
rect 2159 -283 2193 -249
rect 2227 -283 2261 -249
rect 2295 -283 2329 -249
rect 2363 -283 2397 -249
rect 2431 -283 2465 -249
rect 2499 -283 2533 -249
<< poly >>
rect -2500 181 2500 197
rect -2500 147 -2465 181
rect -2431 147 -2397 181
rect -2363 147 -2329 181
rect -2295 147 -2261 181
rect -2227 147 -2193 181
rect -2159 147 -2125 181
rect -2091 147 -2057 181
rect -2023 147 -1989 181
rect -1955 147 -1921 181
rect -1887 147 -1853 181
rect -1819 147 -1785 181
rect -1751 147 -1717 181
rect -1683 147 -1649 181
rect -1615 147 -1581 181
rect -1547 147 -1513 181
rect -1479 147 -1445 181
rect -1411 147 -1377 181
rect -1343 147 -1309 181
rect -1275 147 -1241 181
rect -1207 147 -1173 181
rect -1139 147 -1105 181
rect -1071 147 -1037 181
rect -1003 147 -969 181
rect -935 147 -901 181
rect -867 147 -833 181
rect -799 147 -765 181
rect -731 147 -697 181
rect -663 147 -629 181
rect -595 147 -561 181
rect -527 147 -493 181
rect -459 147 -425 181
rect -391 147 -357 181
rect -323 147 -289 181
rect -255 147 -221 181
rect -187 147 -153 181
rect -119 147 -85 181
rect -51 147 -17 181
rect 17 147 51 181
rect 85 147 119 181
rect 153 147 187 181
rect 221 147 255 181
rect 289 147 323 181
rect 357 147 391 181
rect 425 147 459 181
rect 493 147 527 181
rect 561 147 595 181
rect 629 147 663 181
rect 697 147 731 181
rect 765 147 799 181
rect 833 147 867 181
rect 901 147 935 181
rect 969 147 1003 181
rect 1037 147 1071 181
rect 1105 147 1139 181
rect 1173 147 1207 181
rect 1241 147 1275 181
rect 1309 147 1343 181
rect 1377 147 1411 181
rect 1445 147 1479 181
rect 1513 147 1547 181
rect 1581 147 1615 181
rect 1649 147 1683 181
rect 1717 147 1751 181
rect 1785 147 1819 181
rect 1853 147 1887 181
rect 1921 147 1955 181
rect 1989 147 2023 181
rect 2057 147 2091 181
rect 2125 147 2159 181
rect 2193 147 2227 181
rect 2261 147 2295 181
rect 2329 147 2363 181
rect 2397 147 2431 181
rect 2465 147 2500 181
rect -2500 100 2500 147
rect -2500 -147 2500 -100
rect -2500 -181 -2465 -147
rect -2431 -181 -2397 -147
rect -2363 -181 -2329 -147
rect -2295 -181 -2261 -147
rect -2227 -181 -2193 -147
rect -2159 -181 -2125 -147
rect -2091 -181 -2057 -147
rect -2023 -181 -1989 -147
rect -1955 -181 -1921 -147
rect -1887 -181 -1853 -147
rect -1819 -181 -1785 -147
rect -1751 -181 -1717 -147
rect -1683 -181 -1649 -147
rect -1615 -181 -1581 -147
rect -1547 -181 -1513 -147
rect -1479 -181 -1445 -147
rect -1411 -181 -1377 -147
rect -1343 -181 -1309 -147
rect -1275 -181 -1241 -147
rect -1207 -181 -1173 -147
rect -1139 -181 -1105 -147
rect -1071 -181 -1037 -147
rect -1003 -181 -969 -147
rect -935 -181 -901 -147
rect -867 -181 -833 -147
rect -799 -181 -765 -147
rect -731 -181 -697 -147
rect -663 -181 -629 -147
rect -595 -181 -561 -147
rect -527 -181 -493 -147
rect -459 -181 -425 -147
rect -391 -181 -357 -147
rect -323 -181 -289 -147
rect -255 -181 -221 -147
rect -187 -181 -153 -147
rect -119 -181 -85 -147
rect -51 -181 -17 -147
rect 17 -181 51 -147
rect 85 -181 119 -147
rect 153 -181 187 -147
rect 221 -181 255 -147
rect 289 -181 323 -147
rect 357 -181 391 -147
rect 425 -181 459 -147
rect 493 -181 527 -147
rect 561 -181 595 -147
rect 629 -181 663 -147
rect 697 -181 731 -147
rect 765 -181 799 -147
rect 833 -181 867 -147
rect 901 -181 935 -147
rect 969 -181 1003 -147
rect 1037 -181 1071 -147
rect 1105 -181 1139 -147
rect 1173 -181 1207 -147
rect 1241 -181 1275 -147
rect 1309 -181 1343 -147
rect 1377 -181 1411 -147
rect 1445 -181 1479 -147
rect 1513 -181 1547 -147
rect 1581 -181 1615 -147
rect 1649 -181 1683 -147
rect 1717 -181 1751 -147
rect 1785 -181 1819 -147
rect 1853 -181 1887 -147
rect 1921 -181 1955 -147
rect 1989 -181 2023 -147
rect 2057 -181 2091 -147
rect 2125 -181 2159 -147
rect 2193 -181 2227 -147
rect 2261 -181 2295 -147
rect 2329 -181 2363 -147
rect 2397 -181 2431 -147
rect 2465 -181 2500 -147
rect -2500 -197 2500 -181
<< polycont >>
rect -2465 147 -2431 181
rect -2397 147 -2363 181
rect -2329 147 -2295 181
rect -2261 147 -2227 181
rect -2193 147 -2159 181
rect -2125 147 -2091 181
rect -2057 147 -2023 181
rect -1989 147 -1955 181
rect -1921 147 -1887 181
rect -1853 147 -1819 181
rect -1785 147 -1751 181
rect -1717 147 -1683 181
rect -1649 147 -1615 181
rect -1581 147 -1547 181
rect -1513 147 -1479 181
rect -1445 147 -1411 181
rect -1377 147 -1343 181
rect -1309 147 -1275 181
rect -1241 147 -1207 181
rect -1173 147 -1139 181
rect -1105 147 -1071 181
rect -1037 147 -1003 181
rect -969 147 -935 181
rect -901 147 -867 181
rect -833 147 -799 181
rect -765 147 -731 181
rect -697 147 -663 181
rect -629 147 -595 181
rect -561 147 -527 181
rect -493 147 -459 181
rect -425 147 -391 181
rect -357 147 -323 181
rect -289 147 -255 181
rect -221 147 -187 181
rect -153 147 -119 181
rect -85 147 -51 181
rect -17 147 17 181
rect 51 147 85 181
rect 119 147 153 181
rect 187 147 221 181
rect 255 147 289 181
rect 323 147 357 181
rect 391 147 425 181
rect 459 147 493 181
rect 527 147 561 181
rect 595 147 629 181
rect 663 147 697 181
rect 731 147 765 181
rect 799 147 833 181
rect 867 147 901 181
rect 935 147 969 181
rect 1003 147 1037 181
rect 1071 147 1105 181
rect 1139 147 1173 181
rect 1207 147 1241 181
rect 1275 147 1309 181
rect 1343 147 1377 181
rect 1411 147 1445 181
rect 1479 147 1513 181
rect 1547 147 1581 181
rect 1615 147 1649 181
rect 1683 147 1717 181
rect 1751 147 1785 181
rect 1819 147 1853 181
rect 1887 147 1921 181
rect 1955 147 1989 181
rect 2023 147 2057 181
rect 2091 147 2125 181
rect 2159 147 2193 181
rect 2227 147 2261 181
rect 2295 147 2329 181
rect 2363 147 2397 181
rect 2431 147 2465 181
rect -2465 -181 -2431 -147
rect -2397 -181 -2363 -147
rect -2329 -181 -2295 -147
rect -2261 -181 -2227 -147
rect -2193 -181 -2159 -147
rect -2125 -181 -2091 -147
rect -2057 -181 -2023 -147
rect -1989 -181 -1955 -147
rect -1921 -181 -1887 -147
rect -1853 -181 -1819 -147
rect -1785 -181 -1751 -147
rect -1717 -181 -1683 -147
rect -1649 -181 -1615 -147
rect -1581 -181 -1547 -147
rect -1513 -181 -1479 -147
rect -1445 -181 -1411 -147
rect -1377 -181 -1343 -147
rect -1309 -181 -1275 -147
rect -1241 -181 -1207 -147
rect -1173 -181 -1139 -147
rect -1105 -181 -1071 -147
rect -1037 -181 -1003 -147
rect -969 -181 -935 -147
rect -901 -181 -867 -147
rect -833 -181 -799 -147
rect -765 -181 -731 -147
rect -697 -181 -663 -147
rect -629 -181 -595 -147
rect -561 -181 -527 -147
rect -493 -181 -459 -147
rect -425 -181 -391 -147
rect -357 -181 -323 -147
rect -289 -181 -255 -147
rect -221 -181 -187 -147
rect -153 -181 -119 -147
rect -85 -181 -51 -147
rect -17 -181 17 -147
rect 51 -181 85 -147
rect 119 -181 153 -147
rect 187 -181 221 -147
rect 255 -181 289 -147
rect 323 -181 357 -147
rect 391 -181 425 -147
rect 459 -181 493 -147
rect 527 -181 561 -147
rect 595 -181 629 -147
rect 663 -181 697 -147
rect 731 -181 765 -147
rect 799 -181 833 -147
rect 867 -181 901 -147
rect 935 -181 969 -147
rect 1003 -181 1037 -147
rect 1071 -181 1105 -147
rect 1139 -181 1173 -147
rect 1207 -181 1241 -147
rect 1275 -181 1309 -147
rect 1343 -181 1377 -147
rect 1411 -181 1445 -147
rect 1479 -181 1513 -147
rect 1547 -181 1581 -147
rect 1615 -181 1649 -147
rect 1683 -181 1717 -147
rect 1751 -181 1785 -147
rect 1819 -181 1853 -147
rect 1887 -181 1921 -147
rect 1955 -181 1989 -147
rect 2023 -181 2057 -147
rect 2091 -181 2125 -147
rect 2159 -181 2193 -147
rect 2227 -181 2261 -147
rect 2295 -181 2329 -147
rect 2363 -181 2397 -147
rect 2431 -181 2465 -147
<< locali >>
rect -2660 249 -2533 283
rect -2499 249 -2465 283
rect -2431 249 -2397 283
rect -2363 249 -2329 283
rect -2295 249 -2261 283
rect -2227 249 -2193 283
rect -2159 249 -2125 283
rect -2091 249 -2057 283
rect -2023 249 -1989 283
rect -1955 249 -1921 283
rect -1887 249 -1853 283
rect -1819 249 -1785 283
rect -1751 249 -1717 283
rect -1683 249 -1649 283
rect -1615 249 -1581 283
rect -1547 249 -1513 283
rect -1479 249 -1445 283
rect -1411 249 -1377 283
rect -1343 249 -1309 283
rect -1275 249 -1241 283
rect -1207 249 -1173 283
rect -1139 249 -1105 283
rect -1071 249 -1037 283
rect -1003 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1003 283
rect 1037 249 1071 283
rect 1105 249 1139 283
rect 1173 249 1207 283
rect 1241 249 1275 283
rect 1309 249 1343 283
rect 1377 249 1411 283
rect 1445 249 1479 283
rect 1513 249 1547 283
rect 1581 249 1615 283
rect 1649 249 1683 283
rect 1717 249 1751 283
rect 1785 249 1819 283
rect 1853 249 1887 283
rect 1921 249 1955 283
rect 1989 249 2023 283
rect 2057 249 2091 283
rect 2125 249 2159 283
rect 2193 249 2227 283
rect 2261 249 2295 283
rect 2329 249 2363 283
rect 2397 249 2431 283
rect 2465 249 2499 283
rect 2533 249 2660 283
rect -2660 187 -2626 249
rect 2626 187 2660 249
rect -2660 119 -2626 153
rect -2500 147 -2465 181
rect -2431 147 -2397 181
rect -2359 147 -2329 181
rect -2287 147 -2261 181
rect -2215 147 -2193 181
rect -2143 147 -2125 181
rect -2071 147 -2057 181
rect -1999 147 -1989 181
rect -1927 147 -1921 181
rect -1855 147 -1853 181
rect -1819 147 -1817 181
rect -1751 147 -1745 181
rect -1683 147 -1673 181
rect -1615 147 -1601 181
rect -1547 147 -1529 181
rect -1479 147 -1457 181
rect -1411 147 -1385 181
rect -1343 147 -1313 181
rect -1275 147 -1241 181
rect -1207 147 -1173 181
rect -1135 147 -1105 181
rect -1063 147 -1037 181
rect -991 147 -969 181
rect -919 147 -901 181
rect -847 147 -833 181
rect -775 147 -765 181
rect -703 147 -697 181
rect -631 147 -629 181
rect -595 147 -593 181
rect -527 147 -521 181
rect -459 147 -449 181
rect -391 147 -377 181
rect -323 147 -305 181
rect -255 147 -233 181
rect -187 147 -161 181
rect -119 147 -89 181
rect -51 147 -17 181
rect 17 147 51 181
rect 89 147 119 181
rect 161 147 187 181
rect 233 147 255 181
rect 305 147 323 181
rect 377 147 391 181
rect 449 147 459 181
rect 521 147 527 181
rect 593 147 595 181
rect 629 147 631 181
rect 697 147 703 181
rect 765 147 775 181
rect 833 147 847 181
rect 901 147 919 181
rect 969 147 991 181
rect 1037 147 1063 181
rect 1105 147 1135 181
rect 1173 147 1207 181
rect 1241 147 1275 181
rect 1313 147 1343 181
rect 1385 147 1411 181
rect 1457 147 1479 181
rect 1529 147 1547 181
rect 1601 147 1615 181
rect 1673 147 1683 181
rect 1745 147 1751 181
rect 1817 147 1819 181
rect 1853 147 1855 181
rect 1921 147 1927 181
rect 1989 147 1999 181
rect 2057 147 2071 181
rect 2125 147 2143 181
rect 2193 147 2215 181
rect 2261 147 2287 181
rect 2329 147 2359 181
rect 2397 147 2431 181
rect 2465 147 2500 181
rect 2626 119 2660 153
rect -2660 51 -2626 85
rect -2660 -17 -2626 17
rect -2660 -85 -2626 -51
rect -2546 85 -2512 104
rect -2546 17 -2512 19
rect -2546 -19 -2512 -17
rect -2546 -104 -2512 -85
rect 2512 85 2546 104
rect 2512 17 2546 19
rect 2512 -19 2546 -17
rect 2512 -104 2546 -85
rect 2626 51 2660 85
rect 2626 -17 2660 17
rect 2626 -85 2660 -51
rect -2660 -153 -2626 -119
rect -2500 -181 -2465 -147
rect -2431 -181 -2397 -147
rect -2359 -181 -2329 -147
rect -2287 -181 -2261 -147
rect -2215 -181 -2193 -147
rect -2143 -181 -2125 -147
rect -2071 -181 -2057 -147
rect -1999 -181 -1989 -147
rect -1927 -181 -1921 -147
rect -1855 -181 -1853 -147
rect -1819 -181 -1817 -147
rect -1751 -181 -1745 -147
rect -1683 -181 -1673 -147
rect -1615 -181 -1601 -147
rect -1547 -181 -1529 -147
rect -1479 -181 -1457 -147
rect -1411 -181 -1385 -147
rect -1343 -181 -1313 -147
rect -1275 -181 -1241 -147
rect -1207 -181 -1173 -147
rect -1135 -181 -1105 -147
rect -1063 -181 -1037 -147
rect -991 -181 -969 -147
rect -919 -181 -901 -147
rect -847 -181 -833 -147
rect -775 -181 -765 -147
rect -703 -181 -697 -147
rect -631 -181 -629 -147
rect -595 -181 -593 -147
rect -527 -181 -521 -147
rect -459 -181 -449 -147
rect -391 -181 -377 -147
rect -323 -181 -305 -147
rect -255 -181 -233 -147
rect -187 -181 -161 -147
rect -119 -181 -89 -147
rect -51 -181 -17 -147
rect 17 -181 51 -147
rect 89 -181 119 -147
rect 161 -181 187 -147
rect 233 -181 255 -147
rect 305 -181 323 -147
rect 377 -181 391 -147
rect 449 -181 459 -147
rect 521 -181 527 -147
rect 593 -181 595 -147
rect 629 -181 631 -147
rect 697 -181 703 -147
rect 765 -181 775 -147
rect 833 -181 847 -147
rect 901 -181 919 -147
rect 969 -181 991 -147
rect 1037 -181 1063 -147
rect 1105 -181 1135 -147
rect 1173 -181 1207 -147
rect 1241 -181 1275 -147
rect 1313 -181 1343 -147
rect 1385 -181 1411 -147
rect 1457 -181 1479 -147
rect 1529 -181 1547 -147
rect 1601 -181 1615 -147
rect 1673 -181 1683 -147
rect 1745 -181 1751 -147
rect 1817 -181 1819 -147
rect 1853 -181 1855 -147
rect 1921 -181 1927 -147
rect 1989 -181 1999 -147
rect 2057 -181 2071 -147
rect 2125 -181 2143 -147
rect 2193 -181 2215 -147
rect 2261 -181 2287 -147
rect 2329 -181 2359 -147
rect 2397 -181 2431 -147
rect 2465 -181 2500 -147
rect 2626 -153 2660 -119
rect -2660 -249 -2626 -187
rect 2626 -249 2660 -187
rect -2660 -283 -2533 -249
rect -2499 -283 -2465 -249
rect -2431 -283 -2397 -249
rect -2363 -283 -2329 -249
rect -2295 -283 -2261 -249
rect -2227 -283 -2193 -249
rect -2159 -283 -2125 -249
rect -2091 -283 -2057 -249
rect -2023 -283 -1989 -249
rect -1955 -283 -1921 -249
rect -1887 -283 -1853 -249
rect -1819 -283 -1785 -249
rect -1751 -283 -1717 -249
rect -1683 -283 -1649 -249
rect -1615 -283 -1581 -249
rect -1547 -283 -1513 -249
rect -1479 -283 -1445 -249
rect -1411 -283 -1377 -249
rect -1343 -283 -1309 -249
rect -1275 -283 -1241 -249
rect -1207 -283 -1173 -249
rect -1139 -283 -1105 -249
rect -1071 -283 -1037 -249
rect -1003 -283 -969 -249
rect -935 -283 -901 -249
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
rect 901 -283 935 -249
rect 969 -283 1003 -249
rect 1037 -283 1071 -249
rect 1105 -283 1139 -249
rect 1173 -283 1207 -249
rect 1241 -283 1275 -249
rect 1309 -283 1343 -249
rect 1377 -283 1411 -249
rect 1445 -283 1479 -249
rect 1513 -283 1547 -249
rect 1581 -283 1615 -249
rect 1649 -283 1683 -249
rect 1717 -283 1751 -249
rect 1785 -283 1819 -249
rect 1853 -283 1887 -249
rect 1921 -283 1955 -249
rect 1989 -283 2023 -249
rect 2057 -283 2091 -249
rect 2125 -283 2159 -249
rect 2193 -283 2227 -249
rect 2261 -283 2295 -249
rect 2329 -283 2363 -249
rect 2397 -283 2431 -249
rect 2465 -283 2499 -249
rect 2533 -283 2660 -249
<< viali >>
rect -2465 147 -2431 181
rect -2393 147 -2363 181
rect -2363 147 -2359 181
rect -2321 147 -2295 181
rect -2295 147 -2287 181
rect -2249 147 -2227 181
rect -2227 147 -2215 181
rect -2177 147 -2159 181
rect -2159 147 -2143 181
rect -2105 147 -2091 181
rect -2091 147 -2071 181
rect -2033 147 -2023 181
rect -2023 147 -1999 181
rect -1961 147 -1955 181
rect -1955 147 -1927 181
rect -1889 147 -1887 181
rect -1887 147 -1855 181
rect -1817 147 -1785 181
rect -1785 147 -1783 181
rect -1745 147 -1717 181
rect -1717 147 -1711 181
rect -1673 147 -1649 181
rect -1649 147 -1639 181
rect -1601 147 -1581 181
rect -1581 147 -1567 181
rect -1529 147 -1513 181
rect -1513 147 -1495 181
rect -1457 147 -1445 181
rect -1445 147 -1423 181
rect -1385 147 -1377 181
rect -1377 147 -1351 181
rect -1313 147 -1309 181
rect -1309 147 -1279 181
rect -1241 147 -1207 181
rect -1169 147 -1139 181
rect -1139 147 -1135 181
rect -1097 147 -1071 181
rect -1071 147 -1063 181
rect -1025 147 -1003 181
rect -1003 147 -991 181
rect -953 147 -935 181
rect -935 147 -919 181
rect -881 147 -867 181
rect -867 147 -847 181
rect -809 147 -799 181
rect -799 147 -775 181
rect -737 147 -731 181
rect -731 147 -703 181
rect -665 147 -663 181
rect -663 147 -631 181
rect -593 147 -561 181
rect -561 147 -559 181
rect -521 147 -493 181
rect -493 147 -487 181
rect -449 147 -425 181
rect -425 147 -415 181
rect -377 147 -357 181
rect -357 147 -343 181
rect -305 147 -289 181
rect -289 147 -271 181
rect -233 147 -221 181
rect -221 147 -199 181
rect -161 147 -153 181
rect -153 147 -127 181
rect -89 147 -85 181
rect -85 147 -55 181
rect -17 147 17 181
rect 55 147 85 181
rect 85 147 89 181
rect 127 147 153 181
rect 153 147 161 181
rect 199 147 221 181
rect 221 147 233 181
rect 271 147 289 181
rect 289 147 305 181
rect 343 147 357 181
rect 357 147 377 181
rect 415 147 425 181
rect 425 147 449 181
rect 487 147 493 181
rect 493 147 521 181
rect 559 147 561 181
rect 561 147 593 181
rect 631 147 663 181
rect 663 147 665 181
rect 703 147 731 181
rect 731 147 737 181
rect 775 147 799 181
rect 799 147 809 181
rect 847 147 867 181
rect 867 147 881 181
rect 919 147 935 181
rect 935 147 953 181
rect 991 147 1003 181
rect 1003 147 1025 181
rect 1063 147 1071 181
rect 1071 147 1097 181
rect 1135 147 1139 181
rect 1139 147 1169 181
rect 1207 147 1241 181
rect 1279 147 1309 181
rect 1309 147 1313 181
rect 1351 147 1377 181
rect 1377 147 1385 181
rect 1423 147 1445 181
rect 1445 147 1457 181
rect 1495 147 1513 181
rect 1513 147 1529 181
rect 1567 147 1581 181
rect 1581 147 1601 181
rect 1639 147 1649 181
rect 1649 147 1673 181
rect 1711 147 1717 181
rect 1717 147 1745 181
rect 1783 147 1785 181
rect 1785 147 1817 181
rect 1855 147 1887 181
rect 1887 147 1889 181
rect 1927 147 1955 181
rect 1955 147 1961 181
rect 1999 147 2023 181
rect 2023 147 2033 181
rect 2071 147 2091 181
rect 2091 147 2105 181
rect 2143 147 2159 181
rect 2159 147 2177 181
rect 2215 147 2227 181
rect 2227 147 2249 181
rect 2287 147 2295 181
rect 2295 147 2321 181
rect 2359 147 2363 181
rect 2363 147 2393 181
rect 2431 147 2465 181
rect -2546 51 -2512 53
rect -2546 19 -2512 51
rect -2546 -51 -2512 -19
rect -2546 -53 -2512 -51
rect 2512 51 2546 53
rect 2512 19 2546 51
rect 2512 -51 2546 -19
rect 2512 -53 2546 -51
rect -2465 -181 -2431 -147
rect -2393 -181 -2363 -147
rect -2363 -181 -2359 -147
rect -2321 -181 -2295 -147
rect -2295 -181 -2287 -147
rect -2249 -181 -2227 -147
rect -2227 -181 -2215 -147
rect -2177 -181 -2159 -147
rect -2159 -181 -2143 -147
rect -2105 -181 -2091 -147
rect -2091 -181 -2071 -147
rect -2033 -181 -2023 -147
rect -2023 -181 -1999 -147
rect -1961 -181 -1955 -147
rect -1955 -181 -1927 -147
rect -1889 -181 -1887 -147
rect -1887 -181 -1855 -147
rect -1817 -181 -1785 -147
rect -1785 -181 -1783 -147
rect -1745 -181 -1717 -147
rect -1717 -181 -1711 -147
rect -1673 -181 -1649 -147
rect -1649 -181 -1639 -147
rect -1601 -181 -1581 -147
rect -1581 -181 -1567 -147
rect -1529 -181 -1513 -147
rect -1513 -181 -1495 -147
rect -1457 -181 -1445 -147
rect -1445 -181 -1423 -147
rect -1385 -181 -1377 -147
rect -1377 -181 -1351 -147
rect -1313 -181 -1309 -147
rect -1309 -181 -1279 -147
rect -1241 -181 -1207 -147
rect -1169 -181 -1139 -147
rect -1139 -181 -1135 -147
rect -1097 -181 -1071 -147
rect -1071 -181 -1063 -147
rect -1025 -181 -1003 -147
rect -1003 -181 -991 -147
rect -953 -181 -935 -147
rect -935 -181 -919 -147
rect -881 -181 -867 -147
rect -867 -181 -847 -147
rect -809 -181 -799 -147
rect -799 -181 -775 -147
rect -737 -181 -731 -147
rect -731 -181 -703 -147
rect -665 -181 -663 -147
rect -663 -181 -631 -147
rect -593 -181 -561 -147
rect -561 -181 -559 -147
rect -521 -181 -493 -147
rect -493 -181 -487 -147
rect -449 -181 -425 -147
rect -425 -181 -415 -147
rect -377 -181 -357 -147
rect -357 -181 -343 -147
rect -305 -181 -289 -147
rect -289 -181 -271 -147
rect -233 -181 -221 -147
rect -221 -181 -199 -147
rect -161 -181 -153 -147
rect -153 -181 -127 -147
rect -89 -181 -85 -147
rect -85 -181 -55 -147
rect -17 -181 17 -147
rect 55 -181 85 -147
rect 85 -181 89 -147
rect 127 -181 153 -147
rect 153 -181 161 -147
rect 199 -181 221 -147
rect 221 -181 233 -147
rect 271 -181 289 -147
rect 289 -181 305 -147
rect 343 -181 357 -147
rect 357 -181 377 -147
rect 415 -181 425 -147
rect 425 -181 449 -147
rect 487 -181 493 -147
rect 493 -181 521 -147
rect 559 -181 561 -147
rect 561 -181 593 -147
rect 631 -181 663 -147
rect 663 -181 665 -147
rect 703 -181 731 -147
rect 731 -181 737 -147
rect 775 -181 799 -147
rect 799 -181 809 -147
rect 847 -181 867 -147
rect 867 -181 881 -147
rect 919 -181 935 -147
rect 935 -181 953 -147
rect 991 -181 1003 -147
rect 1003 -181 1025 -147
rect 1063 -181 1071 -147
rect 1071 -181 1097 -147
rect 1135 -181 1139 -147
rect 1139 -181 1169 -147
rect 1207 -181 1241 -147
rect 1279 -181 1309 -147
rect 1309 -181 1313 -147
rect 1351 -181 1377 -147
rect 1377 -181 1385 -147
rect 1423 -181 1445 -147
rect 1445 -181 1457 -147
rect 1495 -181 1513 -147
rect 1513 -181 1529 -147
rect 1567 -181 1581 -147
rect 1581 -181 1601 -147
rect 1639 -181 1649 -147
rect 1649 -181 1673 -147
rect 1711 -181 1717 -147
rect 1717 -181 1745 -147
rect 1783 -181 1785 -147
rect 1785 -181 1817 -147
rect 1855 -181 1887 -147
rect 1887 -181 1889 -147
rect 1927 -181 1955 -147
rect 1955 -181 1961 -147
rect 1999 -181 2023 -147
rect 2023 -181 2033 -147
rect 2071 -181 2091 -147
rect 2091 -181 2105 -147
rect 2143 -181 2159 -147
rect 2159 -181 2177 -147
rect 2215 -181 2227 -147
rect 2227 -181 2249 -147
rect 2287 -181 2295 -147
rect 2295 -181 2321 -147
rect 2359 -181 2363 -147
rect 2363 -181 2393 -147
rect 2431 -181 2465 -147
<< metal1 >>
rect -2496 181 2496 187
rect -2496 147 -2465 181
rect -2431 147 -2393 181
rect -2359 147 -2321 181
rect -2287 147 -2249 181
rect -2215 147 -2177 181
rect -2143 147 -2105 181
rect -2071 147 -2033 181
rect -1999 147 -1961 181
rect -1927 147 -1889 181
rect -1855 147 -1817 181
rect -1783 147 -1745 181
rect -1711 147 -1673 181
rect -1639 147 -1601 181
rect -1567 147 -1529 181
rect -1495 147 -1457 181
rect -1423 147 -1385 181
rect -1351 147 -1313 181
rect -1279 147 -1241 181
rect -1207 147 -1169 181
rect -1135 147 -1097 181
rect -1063 147 -1025 181
rect -991 147 -953 181
rect -919 147 -881 181
rect -847 147 -809 181
rect -775 147 -737 181
rect -703 147 -665 181
rect -631 147 -593 181
rect -559 147 -521 181
rect -487 147 -449 181
rect -415 147 -377 181
rect -343 147 -305 181
rect -271 147 -233 181
rect -199 147 -161 181
rect -127 147 -89 181
rect -55 147 -17 181
rect 17 147 55 181
rect 89 147 127 181
rect 161 147 199 181
rect 233 147 271 181
rect 305 147 343 181
rect 377 147 415 181
rect 449 147 487 181
rect 521 147 559 181
rect 593 147 631 181
rect 665 147 703 181
rect 737 147 775 181
rect 809 147 847 181
rect 881 147 919 181
rect 953 147 991 181
rect 1025 147 1063 181
rect 1097 147 1135 181
rect 1169 147 1207 181
rect 1241 147 1279 181
rect 1313 147 1351 181
rect 1385 147 1423 181
rect 1457 147 1495 181
rect 1529 147 1567 181
rect 1601 147 1639 181
rect 1673 147 1711 181
rect 1745 147 1783 181
rect 1817 147 1855 181
rect 1889 147 1927 181
rect 1961 147 1999 181
rect 2033 147 2071 181
rect 2105 147 2143 181
rect 2177 147 2215 181
rect 2249 147 2287 181
rect 2321 147 2359 181
rect 2393 147 2431 181
rect 2465 147 2496 181
rect -2496 141 2496 147
rect -2552 53 -2506 100
rect -2552 19 -2546 53
rect -2512 19 -2506 53
rect -2552 -19 -2506 19
rect -2552 -53 -2546 -19
rect -2512 -53 -2506 -19
rect -2552 -100 -2506 -53
rect 2506 53 2552 100
rect 2506 19 2512 53
rect 2546 19 2552 53
rect 2506 -19 2552 19
rect 2506 -53 2512 -19
rect 2546 -53 2552 -19
rect 2506 -100 2552 -53
rect -2496 -147 2496 -141
rect -2496 -181 -2465 -147
rect -2431 -181 -2393 -147
rect -2359 -181 -2321 -147
rect -2287 -181 -2249 -147
rect -2215 -181 -2177 -147
rect -2143 -181 -2105 -147
rect -2071 -181 -2033 -147
rect -1999 -181 -1961 -147
rect -1927 -181 -1889 -147
rect -1855 -181 -1817 -147
rect -1783 -181 -1745 -147
rect -1711 -181 -1673 -147
rect -1639 -181 -1601 -147
rect -1567 -181 -1529 -147
rect -1495 -181 -1457 -147
rect -1423 -181 -1385 -147
rect -1351 -181 -1313 -147
rect -1279 -181 -1241 -147
rect -1207 -181 -1169 -147
rect -1135 -181 -1097 -147
rect -1063 -181 -1025 -147
rect -991 -181 -953 -147
rect -919 -181 -881 -147
rect -847 -181 -809 -147
rect -775 -181 -737 -147
rect -703 -181 -665 -147
rect -631 -181 -593 -147
rect -559 -181 -521 -147
rect -487 -181 -449 -147
rect -415 -181 -377 -147
rect -343 -181 -305 -147
rect -271 -181 -233 -147
rect -199 -181 -161 -147
rect -127 -181 -89 -147
rect -55 -181 -17 -147
rect 17 -181 55 -147
rect 89 -181 127 -147
rect 161 -181 199 -147
rect 233 -181 271 -147
rect 305 -181 343 -147
rect 377 -181 415 -147
rect 449 -181 487 -147
rect 521 -181 559 -147
rect 593 -181 631 -147
rect 665 -181 703 -147
rect 737 -181 775 -147
rect 809 -181 847 -147
rect 881 -181 919 -147
rect 953 -181 991 -147
rect 1025 -181 1063 -147
rect 1097 -181 1135 -147
rect 1169 -181 1207 -147
rect 1241 -181 1279 -147
rect 1313 -181 1351 -147
rect 1385 -181 1423 -147
rect 1457 -181 1495 -147
rect 1529 -181 1567 -147
rect 1601 -181 1639 -147
rect 1673 -181 1711 -147
rect 1745 -181 1783 -147
rect 1817 -181 1855 -147
rect 1889 -181 1927 -147
rect 1961 -181 1999 -147
rect 2033 -181 2071 -147
rect 2105 -181 2143 -147
rect 2177 -181 2215 -147
rect 2249 -181 2287 -147
rect 2321 -181 2359 -147
rect 2393 -181 2431 -147
rect 2465 -181 2496 -147
rect -2496 -187 2496 -181
<< properties >>
string FIXED_BBOX -2643 -266 2643 266
<< end >>
