magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -191 2386 191 2472
rect -191 -2386 -105 2386
rect 105 -2386 191 2386
rect -191 -2472 191 -2386
<< psubdiff >>
rect -165 2412 -51 2446
rect -17 2412 17 2446
rect 51 2412 165 2446
rect -165 2329 -131 2412
rect 131 2329 165 2412
rect -165 2261 -131 2295
rect -165 2193 -131 2227
rect -165 2125 -131 2159
rect -165 2057 -131 2091
rect -165 1989 -131 2023
rect -165 1921 -131 1955
rect -165 1853 -131 1887
rect -165 1785 -131 1819
rect -165 1717 -131 1751
rect -165 1649 -131 1683
rect -165 1581 -131 1615
rect -165 1513 -131 1547
rect -165 1445 -131 1479
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect -165 -1479 -131 -1445
rect -165 -1547 -131 -1513
rect -165 -1615 -131 -1581
rect -165 -1683 -131 -1649
rect -165 -1751 -131 -1717
rect -165 -1819 -131 -1785
rect -165 -1887 -131 -1853
rect -165 -1955 -131 -1921
rect -165 -2023 -131 -1989
rect -165 -2091 -131 -2057
rect -165 -2159 -131 -2125
rect -165 -2227 -131 -2193
rect -165 -2295 -131 -2261
rect 131 2261 165 2295
rect 131 2193 165 2227
rect 131 2125 165 2159
rect 131 2057 165 2091
rect 131 1989 165 2023
rect 131 1921 165 1955
rect 131 1853 165 1887
rect 131 1785 165 1819
rect 131 1717 165 1751
rect 131 1649 165 1683
rect 131 1581 165 1615
rect 131 1513 165 1547
rect 131 1445 165 1479
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect 131 -1479 165 -1445
rect 131 -1547 165 -1513
rect 131 -1615 165 -1581
rect 131 -1683 165 -1649
rect 131 -1751 165 -1717
rect 131 -1819 165 -1785
rect 131 -1887 165 -1853
rect 131 -1955 165 -1921
rect 131 -2023 165 -1989
rect 131 -2091 165 -2057
rect 131 -2159 165 -2125
rect 131 -2227 165 -2193
rect 131 -2295 165 -2261
rect -165 -2412 -131 -2329
rect 131 -2412 165 -2329
rect -165 -2446 -51 -2412
rect -17 -2446 17 -2412
rect 51 -2446 165 -2412
<< psubdiffcont >>
rect -51 2412 -17 2446
rect 17 2412 51 2446
rect -165 2295 -131 2329
rect -165 2227 -131 2261
rect -165 2159 -131 2193
rect -165 2091 -131 2125
rect -165 2023 -131 2057
rect -165 1955 -131 1989
rect -165 1887 -131 1921
rect -165 1819 -131 1853
rect -165 1751 -131 1785
rect -165 1683 -131 1717
rect -165 1615 -131 1649
rect -165 1547 -131 1581
rect -165 1479 -131 1513
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect -165 -1513 -131 -1479
rect -165 -1581 -131 -1547
rect -165 -1649 -131 -1615
rect -165 -1717 -131 -1683
rect -165 -1785 -131 -1751
rect -165 -1853 -131 -1819
rect -165 -1921 -131 -1887
rect -165 -1989 -131 -1955
rect -165 -2057 -131 -2023
rect -165 -2125 -131 -2091
rect -165 -2193 -131 -2159
rect -165 -2261 -131 -2227
rect -165 -2329 -131 -2295
rect 131 2295 165 2329
rect 131 2227 165 2261
rect 131 2159 165 2193
rect 131 2091 165 2125
rect 131 2023 165 2057
rect 131 1955 165 1989
rect 131 1887 165 1921
rect 131 1819 165 1853
rect 131 1751 165 1785
rect 131 1683 165 1717
rect 131 1615 165 1649
rect 131 1547 165 1581
rect 131 1479 165 1513
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect 131 -1513 165 -1479
rect 131 -1581 165 -1547
rect 131 -1649 165 -1615
rect 131 -1717 165 -1683
rect 131 -1785 165 -1751
rect 131 -1853 165 -1819
rect 131 -1921 165 -1887
rect 131 -1989 165 -1955
rect 131 -2057 165 -2023
rect 131 -2125 165 -2091
rect 131 -2193 165 -2159
rect 131 -2261 165 -2227
rect 131 -2329 165 -2295
rect -51 -2446 -17 -2412
rect 17 -2446 51 -2412
<< xpolycontact >>
rect -35 1884 35 2316
rect -35 -2316 35 -1884
<< ppolyres >>
rect -35 -1884 35 1884
<< locali >>
rect -165 2412 -51 2446
rect -17 2412 17 2446
rect 51 2412 165 2446
rect -165 2329 -131 2412
rect 131 2329 165 2412
rect -165 2261 -131 2295
rect -165 2193 -131 2227
rect -165 2125 -131 2159
rect -165 2057 -131 2091
rect -165 1989 -131 2023
rect -165 1921 -131 1955
rect -165 1853 -131 1887
rect 131 2261 165 2295
rect 131 2193 165 2227
rect 131 2125 165 2159
rect 131 2057 165 2091
rect 131 1989 165 2023
rect 131 1921 165 1955
rect -165 1785 -131 1819
rect -165 1717 -131 1751
rect -165 1649 -131 1683
rect -165 1581 -131 1615
rect -165 1513 -131 1547
rect -165 1445 -131 1479
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect -165 -1479 -131 -1445
rect -165 -1547 -131 -1513
rect -165 -1615 -131 -1581
rect -165 -1683 -131 -1649
rect -165 -1751 -131 -1717
rect -165 -1819 -131 -1785
rect -165 -1887 -131 -1853
rect 131 1853 165 1887
rect 131 1785 165 1819
rect 131 1717 165 1751
rect 131 1649 165 1683
rect 131 1581 165 1615
rect 131 1513 165 1547
rect 131 1445 165 1479
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect 131 -1479 165 -1445
rect 131 -1547 165 -1513
rect 131 -1615 165 -1581
rect 131 -1683 165 -1649
rect 131 -1751 165 -1717
rect 131 -1819 165 -1785
rect -165 -1955 -131 -1921
rect -165 -2023 -131 -1989
rect -165 -2091 -131 -2057
rect -165 -2159 -131 -2125
rect -165 -2227 -131 -2193
rect -165 -2295 -131 -2261
rect 131 -1887 165 -1853
rect 131 -1955 165 -1921
rect 131 -2023 165 -1989
rect 131 -2091 165 -2057
rect 131 -2159 165 -2125
rect 131 -2227 165 -2193
rect 131 -2295 165 -2261
rect -165 -2412 -131 -2329
rect 131 -2412 165 -2329
rect -165 -2446 -51 -2412
rect -17 -2446 17 -2412
rect 51 -2446 165 -2412
<< viali >>
rect -17 2262 17 2296
rect -17 2190 17 2224
rect -17 2118 17 2152
rect -17 2046 17 2080
rect -17 1974 17 2008
rect -17 1902 17 1936
rect -17 -1937 17 -1903
rect -17 -2009 17 -1975
rect -17 -2081 17 -2047
rect -17 -2153 17 -2119
rect -17 -2225 17 -2191
rect -17 -2297 17 -2263
<< metal1 >>
rect -25 2296 25 2310
rect -25 2262 -17 2296
rect 17 2262 25 2296
rect -25 2224 25 2262
rect -25 2190 -17 2224
rect 17 2190 25 2224
rect -25 2152 25 2190
rect -25 2118 -17 2152
rect 17 2118 25 2152
rect -25 2080 25 2118
rect -25 2046 -17 2080
rect 17 2046 25 2080
rect -25 2008 25 2046
rect -25 1974 -17 2008
rect 17 1974 25 2008
rect -25 1936 25 1974
rect -25 1902 -17 1936
rect 17 1902 25 1936
rect -25 1889 25 1902
rect -25 -1903 25 -1889
rect -25 -1937 -17 -1903
rect 17 -1937 25 -1903
rect -25 -1975 25 -1937
rect -25 -2009 -17 -1975
rect 17 -2009 25 -1975
rect -25 -2047 25 -2009
rect -25 -2081 -17 -2047
rect 17 -2081 25 -2047
rect -25 -2119 25 -2081
rect -25 -2153 -17 -2119
rect 17 -2153 25 -2119
rect -25 -2191 25 -2153
rect -25 -2225 -17 -2191
rect 17 -2225 25 -2191
rect -25 -2263 25 -2225
rect -25 -2297 -17 -2263
rect 17 -2297 25 -2263
rect -25 -2310 25 -2297
<< properties >>
string FIXED_BBOX -148 -2429 148 2429
<< end >>
