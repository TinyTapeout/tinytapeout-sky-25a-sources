magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 576 240
<< ptap >>
rect -48 60 624 100
rect -48 100 624 140
rect -48 140 624 180
rect -48 180 48 220
rect 528 180 624 220
rect -48 220 48 260
rect 528 220 624 260
<< locali >>
rect -48 60 624 100
rect -48 100 624 140
rect -48 140 624 180
rect -48 180 48 220
rect 528 180 624 220
rect -48 220 48 260
rect 528 220 624 260
<< ptapc >>
rect 80 100 464 140
<< pwell >>
rect -92 -64 668 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 576 240
<< end >>
