magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 1024 1280
use JNWATR_PCH_2CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 512 240
use JNWATR_PCH_2C1F2 xa2 
transform 1 0 0 0 1 240
box 0 240 512 640
use JNWATR_PCH_2C5F0 xa3 
transform 1 0 0 0 1 640
box 0 640 512 1040
use JNWATR_PCH_2CTAPTOP xa4 
transform 1 0 0 0 1 1040
box 0 1040 512 1280
use JNWATR_PCH_2CTAPBOT xb1 
transform 1 0 512 0 1 0
box 512 0 1024 240
use JNWATR_PCH_2C1F2 xb2 
transform 1 0 512 0 1 240
box 512 240 1024 640
use JNWATR_PCH_2C5F0 xb3 
transform 1 0 512 0 1 640
box 512 640 1024 1040
use JNWATR_PCH_2CTAPTOP xb4 
transform 1 0 512 0 1 1040
box 512 1040 1024 1280
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1024 1280
<< end >>
