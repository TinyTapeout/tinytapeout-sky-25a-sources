magic
tech sky130A
magscale 1 1
timestamp 1737500400
<< checkpaint >>
rect 0 0 88 88
<< locali >>
rect 0 0 84 84
<< viali >>
rect 6 6 32 32
rect 6 52 32 78
rect 52 6 78 32
rect 52 52 78 78
<< m1 >>
rect 0 0 88 88
<< v1 >>
rect 6 6 34 34
rect 6 54 34 82
rect 54 6 82 34
rect 54 54 82 82
<< m2 >>
rect 0 0 88 88
<< v2 >>
rect 6 6 34 34
rect 6 54 34 82
rect 54 6 82 34
rect 54 54 82 82
<< m3 >>
rect 0 0 88 88
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 88 88
<< end >>
