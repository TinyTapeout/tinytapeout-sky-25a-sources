magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 1408 1280
use JNWATR_NCH_8CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 704 240
use JNWATR_NCH_8C1F2 xa2 
transform 1 0 0 0 1 240
box 0 240 704 640
use JNWATR_NCH_8C5F0 xa3 
transform 1 0 0 0 1 640
box 0 640 704 1040
use JNWATR_NCH_8CTAPTOP xa4 
transform 1 0 0 0 1 1040
box 0 1040 704 1280
use JNWATR_NCH_8CTAPBOT xb1 
transform 1 0 704 0 1 0
box 704 0 1408 240
use JNWATR_NCH_8C1F2 xb2 
transform 1 0 704 0 1 240
box 704 240 1408 640
use JNWATR_NCH_8C5F0 xb3 
transform 1 0 704 0 1 640
box 704 640 1408 1040
use JNWATR_NCH_8CTAPTOP xb4 
transform 1 0 704 0 1 1040
box 704 1040 1408 1280
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1408 1280
<< end >>
