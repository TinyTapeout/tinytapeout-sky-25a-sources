magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 832 240
<< ptap >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 784 20 880 60
rect -48 60 880 100
rect -48 100 880 140
rect -48 140 880 180
<< locali >>
rect -48 -20 48 20
rect 784 -20 880 20
rect -48 20 48 60
rect 784 20 880 60
rect -48 60 880 100
rect -48 100 880 140
rect -48 140 880 180
<< ptapc >>
rect 80 100 752 140
<< pwell >>
rect -92 -64 924 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 832 240
<< end >>
