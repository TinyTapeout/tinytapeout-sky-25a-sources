magic
tech sky130A
magscale 1 2
timestamp 1757256347
<< nwell >>
rect -308 -362 308 362
<< mvpmos >>
rect -50 -64 50 136
<< mvpdiff >>
rect -108 124 -50 136
rect -108 -52 -96 124
rect -62 -52 -50 124
rect -108 -64 -50 -52
rect 50 124 108 136
rect 50 -52 62 124
rect 96 -52 108 124
rect 50 -64 108 -52
<< mvpdiffc >>
rect -96 -52 -62 124
rect 62 -52 96 124
<< mvnsubdiff >>
rect -242 284 242 296
rect -242 250 -134 284
rect 134 250 242 284
rect -242 238 242 250
rect -242 188 -184 238
rect -242 -188 -230 188
rect -196 -188 -184 188
rect 184 188 242 238
rect -242 -238 -184 -188
rect 184 -188 196 188
rect 230 -188 242 188
rect 184 -238 242 -188
rect -242 -250 242 -238
rect -242 -284 -134 -250
rect 134 -284 242 -250
rect -242 -296 242 -284
<< mvnsubdiffcont >>
rect -134 250 134 284
rect -230 -188 -196 188
rect 196 -188 230 188
rect -134 -284 134 -250
<< poly >>
rect -50 136 50 162
rect -50 -111 50 -64
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect -50 -161 50 -145
<< polycont >>
rect -34 -145 34 -111
<< locali >>
rect -230 250 -134 284
rect 134 250 230 284
rect -230 188 -196 250
rect 196 188 230 250
rect -96 124 -62 140
rect -96 -68 -62 -52
rect 62 124 96 140
rect 62 -68 96 -52
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect -230 -250 -196 -188
rect 196 -250 230 -188
rect -230 -284 -134 -250
rect 134 -284 230 -250
<< viali >>
rect -96 -52 -62 124
rect 62 -52 96 124
rect -34 -145 34 -111
<< metal1 >>
rect -102 124 -56 136
rect -102 -52 -96 124
rect -62 -52 -56 124
rect -102 -64 -56 -52
rect 56 124 102 136
rect 56 -52 62 124
rect 96 -52 102 124
rect 56 -64 102 -52
rect -46 -111 46 -105
rect -46 -145 -34 -111
rect 34 -145 46 -111
rect -46 -151 46 -145
<< labels >>
rlabel mvnsubdiffcont 0 -267 0 -267 0 B
port 1 nsew
rlabel mvpdiffc -79 36 -79 36 0 D
port 2 nsew
rlabel mvpdiffc 79 36 79 36 0 S
port 3 nsew
rlabel polycont 0 -128 0 -128 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -213 -267 213 267
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
