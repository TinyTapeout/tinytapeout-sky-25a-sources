** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tt_um_13hihi31_tdc.sch
.subckt tt_um_13hihi31_tdc clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
*.PININFO VDPWR:B ua[0]:I uo_out[0]:O VGND:B ui_in[0]:I uo_out[1]:O uo_out[2]:O uo_out[3]:O uo_out[4]:O uo_out[5]:O uo_out[6]:O
*+ uo_out[7]:O ui_in[1]:I ui_in[2]:I ui_in[3]:I ui_in[4]:I ui_in[5]:I ui_in[6]:I ui_in[7]:I uio_in[0]:I uio_in[1]:I uio_in[2]:I uio_in[3]:I
*+ uio_in[4]:I uio_in[5]:I uio_in[6]:I uio_in[7]:I uio_out[0]:O uio_out[1]:O uio_out[2]:O uio_out[3]:O uio_out[4]:O uio_out[5]:O uio_out[6]:O
*+ uio_out[7]:O uio_oe[0]:O uio_oe[1]:O uio_oe[2]:O uio_oe[3]:O uio_oe[4]:O uio_oe[5]:O uio_oe[6]:O uio_oe[7]:O ua[1]:I ua[2]:I ua[3]:I ua[4]:I
*+ ua[5]:I ua[6]:I ua[7]:I ena:I clk:I rst_n:I
x2 ua[0] uio_in[5] uio_in[1] uio_in[2] uio_in[3] uio_in[4] start VDPWR VGND input_stage
x4 stop uio_in[0] ui_in[7] ui_in[6] ui_in[5] ui_in[4] stop_delayed VDPWR VGND variable_delay_short
x6 start start_delayed VDPWR VGND variable_delay_dummy
x1 ua[0] VDPWR ui_in[0] ui_in[1] ui_in[2] ui_in[3] stop VDPWR VGND input_stage
x3 start_delayed stop_delayed uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
+ tdc_vernier_buffers
* noconn uio_out[0]
* noconn uio_out[1]
* noconn uio_out[2]
* noconn uio_out[3]
* noconn uio_out[4]
* noconn uio_out[5]
* noconn uio_out[6]
* noconn uio_out[7]
* noconn uio_oe[0]
* noconn uio_oe[1]
* noconn uio_oe[2]
* noconn uio_oe[3]
* noconn uio_oe[4]
* noconn uio_oe[5]
* noconn uio_oe[6]
* noconn uio_oe[7]
* noconn uio_in[7]
* noconn uio_in[6]
* noconn ua[7]
* noconn ua[6]
* noconn ua[5]
* noconn ua[4]
* noconn ua[3]
* noconn ua[2]
* noconn ua[1]
* noconn rst_n
* noconn clk
* noconn ena
.ends

* expanding   symbol:  input_stage.sym # of pins=9
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/input_stage.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/input_stage.sch
.subckt input_stage in en t0 t1 t2 t3 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B t0:I t1:I t2:I t3:I en:I
x1 en in net1 VDD VSS nand_gate
x2 net1 net2 VDD VSS inverter_2
x3 net2 t0 t1 net3 VDD VSS fine_delay
x4 net3 t2 t3 out VDD VSS fine_delay
.ends


* expanding   symbol:  variable_delay_short.sym # of pins=9
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_short.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_short.sch
.subckt variable_delay_short in en_0 en_1 en_2 en_3 en_4 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en_0:I en_1:I en_2:I en_3:I en_4:I
x1 in en_0 out_1 forward_0 out VDD VSS variable_delay_unit
x2 forward_0 en_1 out_2 forward_1 out_1 VDD VSS variable_delay_unit
x3 forward_1 en_2 out_3 forward_2 out_2 VDD VSS variable_delay_unit
x4 forward_2 en_3 out_4 forward_3 out_3 VDD VSS variable_delay_unit
x9 forward_4 VDD VSS net1 out_5 VDD VSS variable_delay_unit
x5 forward_3 en_4 out_5 forward_4 out_4 VDD VSS variable_delay_unit
.ends


* expanding   symbol:  variable_delay_dummy.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_dummy.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_dummy.sch
.subckt variable_delay_dummy in out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B
x1 in VDD out_1 forward_0 out VDD VSS variable_delay_unit
x9 forward_0 VDD VSS net1 out_1 VDD VSS variable_delay_unit
.ends


* expanding   symbol:  tdc_vernier_buffers.sym # of pins=12
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tdc_vernier_buffers.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tdc_vernier_buffers.sch
.subckt tdc_vernier_buffers start stop term_0 term_1 term_2 term_3 term_4 term_5 term_6 term_7 VDD VSS
*.PININFO VDD:B VSS:B start:I stop:I term_0:O term_1:O term_2:O term_3:O term_4:O term_5:O term_6:O term_7:O
x3 start_delay start_buff start_pos start_neg VDD VSS diff_gen
x19 start_pos start_neg stop_strong term_0 term_1 term_2 term_3 term_4 term_5 term_6 term_7 VDD VSS vernier_delay_line
x1 stop stop_strong VDD VSS stop_buffer
x2 start start_delay start_buff VDD VSS start_buffer
.ends


* expanding   symbol:  nand_gate.sym # of pins=5
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/nand_gate.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/nand_gate.sch
.subckt nand_gate a b out VDD VSS
*.PININFO VDD:B a:I out:O VSS:B b:I
XM7 out a net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 out a VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net1 b VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 out b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
.ends


* expanding   symbol:  inverter_2.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sch
.subckt inverter_2 in out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  fine_delay.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/fine_delay.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/fine_delay.sch
.subckt fine_delay in t0 t1 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B t0:I t1:I
XM1 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net3 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net3 t1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM8 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM9 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net2 in net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net2 t0 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  variable_delay_unit.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_unit.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_unit.sch
.subckt variable_delay_unit in en back forward out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en:I back:I forward:O
x1 forward en nen out VDD VSS tristate_inverter
x2 in forward VDD VSS inverter_2
x3 en nen VDD VSS inverter_2
x4 back nen en out VDD VSS tristate_inverter
.ends


* expanding   symbol:  diff_gen.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/diff_gen.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/diff_gen.sch
.subckt diff_gen in_delay in_buff out_pos out_neg VDD VSS
*.PININFO VDD:B VSS:B in_delay:I out_pos:O in_buff:I out_neg:O
x1 out_1_1 in_buff in_delay VDD out_2_1 VSS delay_unit
x2 out_1_2 out_1_1 out_2_1 VDD out_2_2 VSS delay_unit
x3 out_1_3 out_1_2 out_2_2 VDD out_2_3 VSS delay_unit
x4 out_1_4 out_1_3 out_2_3 VDD out_2_4 VSS delay_unit
x5 out_1_5 out_1_4 out_2_4 VDD out_2_5 VSS delay_unit
x6 out_1_6 out_1_5 out_2_5 VDD out_2_6 VSS delay_unit
x7 out_pos out_1_6 out_2_6 VDD out_neg VSS delay_unit
.ends


* expanding   symbol:  vernier_delay_line.sym # of pins=13
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/vernier_delay_line.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/vernier_delay_line.sch
.subckt vernier_delay_line start_pos start_neg stop_strong term_0 term_1 term_2 term_3 term_4 term_5 term_6 term_7 VDD VSS
*.PININFO VDD:B VSS:B start_pos:I stop_strong:I term_0:O term_1:O term_2:O term_3:O term_4:O term_5:O term_6:O term_7:O
*+ start_neg:I
x1 delay_pos_0 start_pos start_neg VDD delay_neg_0 VSS delay_unit
x2 delay_pos_0 delay_neg_0 stop_strong term_0 net1 VDD VSS saff
x4 delay_pos_1 delay_neg_1 stop_strong term_1 net2 VDD VSS saff
x5 delay_pos_1 delay_pos_0 delay_neg_0 VDD delay_neg_1 VSS delay_unit
x6 delay_pos_2 delay_pos_1 delay_neg_1 VDD delay_neg_2 VSS delay_unit
x7 delay_pos_3 delay_pos_2 delay_neg_2 VDD delay_neg_3 VSS delay_unit
x8 delay_pos_2 delay_neg_2 stop_strong term_2 net3 VDD VSS saff
x9 delay_pos_4 delay_pos_3 delay_neg_3 VDD delay_neg_4 VSS delay_unit
x10 delay_pos_3 delay_neg_3 stop_strong term_3 net4 VDD VSS saff
x11 delay_pos_4 delay_neg_4 stop_strong term_4 net5 VDD VSS saff
x12 delay_pos_5 delay_pos_4 delay_neg_4 VDD delay_neg_5 VSS delay_unit
x13 delay_pos_5 delay_neg_5 stop_strong term_5 net6 VDD VSS saff
x14 delay_pos_6 delay_pos_5 delay_neg_5 VDD delay_neg_6 VSS delay_unit
x15 delay_pos_6 delay_neg_6 stop_strong term_6 net7 VDD VSS saff
x16 delay_pos_7 delay_pos_6 delay_neg_6 VDD delay_neg_7 VSS delay_unit
x17 delay_pos_7 delay_neg_7 stop_strong term_7 net8 VDD VSS saff
x18 net9 delay_pos_7 delay_neg_7 VDD net10 VSS delay_unit
.ends


* expanding   symbol:  stop_buffer.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/stop_buffer.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/stop_buffer.sch
.subckt stop_buffer stop stop_strong VDD VSS
*.PININFO VDD:B VSS:B stop:I stop_strong:O
XM7 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM8 net1 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 net3 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM10 net3 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net4 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM12 net4 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 net5 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM14 net5 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM15 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM16 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM17 net7 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM18 net7 net6 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM19 net8 net7 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=12 nf=1 m=1
XM20 net8 net7 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 m=1
XM21 stop_strong net8 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=48 nf=1 m=1
XM22 stop_strong net8 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=1 m=1
XM23 net9 stop VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM24 net9 stop VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM25 net2 net9 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM26 net2 net9 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  start_buffer.sym # of pins=5
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/start_buffer.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/start_buffer.sch
.subckt start_buffer start start_delay start_buff VDD VSS
*.PININFO VDD:B VSS:B start:I start_delay:O start_buff:O
XM1 net1 start VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net1 start VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 start_buff net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=12 nf=1 m=1
XM4 start_buff net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 m=1
XM5 start_delay start_buff VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM6 start_delay start_buff VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
.ends


* expanding   symbol:  tristate_inverter.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tristate_inverter.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tristate_inverter.sch
.subckt tristate_inverter in en nen out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en:I nen:I
XM5 out in net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM7 out in net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 net2 nen VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM2 net1 en VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
.ends


* expanding   symbol:  delay_unit.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/delay_unit.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/delay_unit.sch
.subckt delay_unit out_1 in_1 in_2 VDD out_2 VSS
*.PININFO VDD:B in_1:I out_1:O VSS:B in_2:I out_2:O
XM5 out_2 in_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM7 out_2 in_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM1 out_1 in_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM2 out_1 in_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM3 in_1 in_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM4 in_1 in_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 in_2 in_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM8 in_2 in_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  saff.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/saff.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/saff.sch
.subckt saff d nd clk q nq VDD VSS
*.PININFO VDD:B d:I q:O VSS:B nd:I clk:I nq:O
XM2 net3 q VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 left_latch_1 clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM4 right_latch_1 clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM5 right_latch_1 left_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM6 left_latch_1 right_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM7 right_latch_1 left_latch_1 net7 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=6 nf=2 m=1
XM8 left_latch_1 right_latch_1 net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=6 nf=2 m=1
XM9 net6 clk VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=15 nf=3 m=1
XM10 net7 nd net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=12 nf=3 m=1
XM11 net5 d net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=12 nf=3 m=1
XM12 right_latch_2 left_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM13 right_latch_2 left_latch_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 left_latch_2 right_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM15 left_latch_2 right_latch_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM16 q left_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM17 q left_latch_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM18 nq right_latch_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM19 nq right_latch_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM20 net2 q VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM21 nq right_latch_2 net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM22 q left_latch_2 net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM23 net1 nq VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM24 q left_latch_1 net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM25 nq right_latch_1 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM26 net4 nq VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
