magic
tech sky130A
magscale 1 2
timestamp 1752183586
<< nwell >>
rect -60 -40 780 270
<< pwell >>
rect -40 -302 760 -88
<< nmos >>
rect 50 -250 80 -126
rect 250 -250 280 -126
rect 346 -250 376 -126
rect 546 -250 576 -126
rect 650 -250 680 -126
<< pmos >>
rect 50 0 80 190
rect 250 0 280 190
rect 450 0 480 190
rect 650 0 680 190
<< ndiff >>
rect -8 -150 50 -126
rect -8 -230 0 -150
rect 34 -230 50 -150
rect -8 -250 50 -230
rect 80 -140 138 -126
rect 80 -220 96 -140
rect 130 -220 138 -140
rect 80 -250 138 -220
rect 192 -160 250 -126
rect 192 -220 200 -160
rect 234 -220 250 -160
rect 192 -250 250 -220
rect 280 -180 346 -126
rect 280 -220 296 -180
rect 330 -220 346 -180
rect 280 -250 346 -220
rect 376 -160 434 -126
rect 376 -230 392 -160
rect 426 -230 434 -160
rect 376 -250 434 -230
rect 488 -160 546 -126
rect 488 -220 496 -160
rect 530 -220 546 -160
rect 488 -250 546 -220
rect 576 -206 650 -126
rect 576 -240 596 -206
rect 634 -240 650 -206
rect 576 -250 650 -240
rect 680 -160 738 -126
rect 680 -220 696 -160
rect 730 -220 738 -160
rect 680 -250 738 -220
<< pdiff >>
rect -8 160 50 190
rect -8 40 0 160
rect 34 40 50 160
rect -8 0 50 40
rect 80 160 138 190
rect 80 40 96 160
rect 130 40 138 160
rect 80 0 138 40
rect 192 160 250 190
rect 192 100 200 160
rect 234 100 250 160
rect 192 0 250 100
rect 280 160 338 190
rect 280 100 296 160
rect 330 100 338 160
rect 280 0 338 100
rect 392 160 450 190
rect 392 40 400 160
rect 434 40 450 160
rect 392 0 450 40
rect 480 160 538 190
rect 480 40 496 160
rect 530 40 538 160
rect 480 0 538 40
rect 592 160 650 190
rect 592 100 600 160
rect 634 100 650 160
rect 592 0 650 100
rect 680 160 738 190
rect 680 100 696 160
rect 730 100 738 160
rect 680 0 738 100
<< ndiffc >>
rect 0 -230 34 -150
rect 96 -220 130 -140
rect 200 -220 234 -160
rect 296 -220 330 -180
rect 392 -230 426 -160
rect 496 -220 530 -160
rect 596 -240 634 -206
rect 696 -220 730 -160
<< pdiffc >>
rect 0 40 34 160
rect 96 40 130 160
rect 200 100 234 160
rect 296 100 330 160
rect 400 40 434 160
rect 496 40 530 160
rect 600 100 634 160
rect 696 100 730 160
<< poly >>
rect 50 190 80 216
rect 250 190 280 216
rect 450 190 480 218
rect 650 190 680 216
rect 50 -28 80 0
rect 250 -28 280 0
rect 450 -28 480 0
rect 50 -48 280 -28
rect 50 -82 170 -48
rect 230 -82 280 -48
rect 50 -102 280 -82
rect 50 -126 80 -102
rect 250 -126 280 -102
rect 346 -48 576 -28
rect 346 -82 370 -48
rect 430 -82 576 -48
rect 346 -102 576 -82
rect 346 -126 376 -102
rect 546 -126 576 -102
rect 650 -38 680 0
rect 650 -48 724 -38
rect 650 -82 670 -48
rect 704 -82 724 -48
rect 650 -92 724 -82
rect 650 -126 680 -92
rect 50 -278 80 -250
rect 250 -278 280 -250
rect 346 -278 376 -250
rect 546 -278 576 -250
rect 650 -278 680 -250
<< polycont >>
rect 170 -82 230 -48
rect 370 -82 430 -48
rect 670 -82 704 -48
<< locali >>
rect 0 160 34 180
rect 0 20 34 40
rect 96 160 130 180
rect 200 160 234 180
rect 296 160 330 180
rect 296 80 330 100
rect 400 160 434 260
rect 96 36 130 40
rect 96 2 350 36
rect 400 20 434 40
rect 496 160 530 180
rect 596 160 634 180
rect 596 80 634 100
rect 696 160 730 180
rect 696 80 730 100
rect 0 -150 34 -130
rect 0 -250 34 -230
rect 96 -140 130 2
rect 316 -32 350 2
rect 496 4 530 40
rect 496 -30 684 4
rect 164 -48 236 -32
rect 230 -82 236 -48
rect 164 -98 236 -82
rect 316 -48 450 -32
rect 316 -82 370 -48
rect 430 -64 450 -48
rect 650 -42 684 -30
rect 650 -48 724 -42
rect 430 -82 616 -64
rect 316 -98 616 -82
rect 650 -82 670 -48
rect 704 -82 724 -48
rect 650 -88 724 -82
rect 582 -122 616 -98
rect 96 -240 130 -220
rect 200 -160 234 -140
rect 392 -160 426 -140
rect 200 -240 234 -220
rect 296 -180 330 -160
rect 392 -250 426 -230
rect 496 -160 530 -140
rect 582 -156 730 -122
rect 696 -160 730 -156
rect 496 -240 530 -220
rect 696 -240 730 -220
rect 596 -256 634 -240
<< viali >>
rect 0 40 34 160
rect 200 100 234 140
rect 200 80 234 100
rect 296 100 330 160
rect 400 40 434 120
rect 496 40 530 120
rect 596 100 600 160
rect 600 100 634 160
rect 696 100 730 160
rect 0 -230 34 -150
rect 164 -82 170 -48
rect 170 -82 198 -48
rect 200 -220 234 -160
rect 296 -220 330 -200
rect 296 -240 330 -220
rect 392 -230 426 -160
rect 496 -220 530 -160
rect 596 -206 634 -190
rect 596 -240 634 -206
<< metal1 >>
rect -40 194 40 274
rect -6 160 40 194
rect 290 170 640 210
rect 290 160 336 170
rect -6 40 0 160
rect 34 40 40 160
rect -6 28 40 40
rect 194 140 240 160
rect 194 80 200 140
rect 234 80 240 140
rect 290 100 296 160
rect 330 100 336 160
rect 590 160 640 170
rect 290 88 336 100
rect 394 120 440 140
rect 194 64 240 80
rect 246 12 266 64
rect 194 0 266 12
rect 394 40 400 120
rect 434 40 440 120
rect 394 0 440 40
rect 130 -42 204 -36
rect 130 -94 142 -42
rect 194 -48 204 -42
rect 198 -82 204 -48
rect 194 -94 204 -82
rect -6 -150 100 -138
rect -6 -230 0 -150
rect 34 -170 100 -150
rect 34 -230 40 -170
rect 92 -230 100 -170
rect -6 -254 100 -230
rect -40 -334 100 -254
rect 130 -280 164 -94
rect 232 -124 266 0
rect 194 -160 266 -124
rect 294 -40 440 0
rect 490 120 542 140
rect 490 64 496 120
rect 530 64 542 120
rect 194 -220 200 -160
rect 234 -220 240 -160
rect 294 -188 336 -40
rect 194 -240 240 -220
rect 290 -200 336 -188
rect 290 -240 296 -200
rect 330 -240 336 -200
rect 290 -252 336 -240
rect 386 -160 438 -148
rect 386 -170 392 -160
rect 426 -170 438 -160
rect 386 -242 438 -230
rect 490 -160 542 12
rect 490 -220 496 -160
rect 530 -220 542 -160
rect 490 -240 542 -220
rect 590 100 596 160
rect 634 100 640 160
rect 590 -190 640 100
rect 684 160 736 172
rect 684 100 696 160
rect 730 100 736 160
rect 684 -42 736 100
rect 684 -106 736 -94
rect 590 -240 596 -190
rect 634 -240 640 -190
rect 590 -252 640 -240
rect 130 -310 336 -280
<< via1 >>
rect 194 12 246 64
rect 142 -48 194 -42
rect 142 -82 164 -48
rect 164 -82 194 -48
rect 142 -94 194 -82
rect 40 -230 92 -170
rect 490 40 496 64
rect 496 40 530 64
rect 530 40 542 64
rect 490 12 542 40
rect 386 -230 392 -170
rect 392 -230 426 -170
rect 426 -230 438 -170
rect 684 -94 736 -42
<< metal2 >>
rect 194 64 542 76
rect 246 12 490 64
rect 194 0 542 12
rect 130 -94 142 -42
rect 194 -94 684 -42
rect 736 -94 742 -42
rect 40 -170 438 -150
rect 92 -230 386 -170
rect 40 -250 438 -230
<< properties >>
string MASKHINTS_PSDM -33 0 763 280
<< end >>
