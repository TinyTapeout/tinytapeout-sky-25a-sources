magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -77 981 -19 987
rect 115 981 173 987
rect -77 947 -65 981
rect 115 947 127 981
rect -77 941 -19 947
rect 115 941 173 947
rect -173 -947 -115 -941
rect 19 -947 77 -941
rect -173 -981 -161 -947
rect 19 -981 31 -947
rect -173 -987 -115 -981
rect 19 -987 77 -981
<< nwell >>
rect -359 -1119 359 1119
<< pmos >>
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
<< pdiff >>
rect -221 867 -159 900
rect -221 833 -209 867
rect -175 833 -159 867
rect -221 799 -159 833
rect -221 765 -209 799
rect -175 765 -159 799
rect -221 731 -159 765
rect -221 697 -209 731
rect -175 697 -159 731
rect -221 663 -159 697
rect -221 629 -209 663
rect -175 629 -159 663
rect -221 595 -159 629
rect -221 561 -209 595
rect -175 561 -159 595
rect -221 527 -159 561
rect -221 493 -209 527
rect -175 493 -159 527
rect -221 459 -159 493
rect -221 425 -209 459
rect -175 425 -159 459
rect -221 391 -159 425
rect -221 357 -209 391
rect -175 357 -159 391
rect -221 323 -159 357
rect -221 289 -209 323
rect -175 289 -159 323
rect -221 255 -159 289
rect -221 221 -209 255
rect -175 221 -159 255
rect -221 187 -159 221
rect -221 153 -209 187
rect -175 153 -159 187
rect -221 119 -159 153
rect -221 85 -209 119
rect -175 85 -159 119
rect -221 51 -159 85
rect -221 17 -209 51
rect -175 17 -159 51
rect -221 -17 -159 17
rect -221 -51 -209 -17
rect -175 -51 -159 -17
rect -221 -85 -159 -51
rect -221 -119 -209 -85
rect -175 -119 -159 -85
rect -221 -153 -159 -119
rect -221 -187 -209 -153
rect -175 -187 -159 -153
rect -221 -221 -159 -187
rect -221 -255 -209 -221
rect -175 -255 -159 -221
rect -221 -289 -159 -255
rect -221 -323 -209 -289
rect -175 -323 -159 -289
rect -221 -357 -159 -323
rect -221 -391 -209 -357
rect -175 -391 -159 -357
rect -221 -425 -159 -391
rect -221 -459 -209 -425
rect -175 -459 -159 -425
rect -221 -493 -159 -459
rect -221 -527 -209 -493
rect -175 -527 -159 -493
rect -221 -561 -159 -527
rect -221 -595 -209 -561
rect -175 -595 -159 -561
rect -221 -629 -159 -595
rect -221 -663 -209 -629
rect -175 -663 -159 -629
rect -221 -697 -159 -663
rect -221 -731 -209 -697
rect -175 -731 -159 -697
rect -221 -765 -159 -731
rect -221 -799 -209 -765
rect -175 -799 -159 -765
rect -221 -833 -159 -799
rect -221 -867 -209 -833
rect -175 -867 -159 -833
rect -221 -900 -159 -867
rect -129 867 -63 900
rect -129 833 -113 867
rect -79 833 -63 867
rect -129 799 -63 833
rect -129 765 -113 799
rect -79 765 -63 799
rect -129 731 -63 765
rect -129 697 -113 731
rect -79 697 -63 731
rect -129 663 -63 697
rect -129 629 -113 663
rect -79 629 -63 663
rect -129 595 -63 629
rect -129 561 -113 595
rect -79 561 -63 595
rect -129 527 -63 561
rect -129 493 -113 527
rect -79 493 -63 527
rect -129 459 -63 493
rect -129 425 -113 459
rect -79 425 -63 459
rect -129 391 -63 425
rect -129 357 -113 391
rect -79 357 -63 391
rect -129 323 -63 357
rect -129 289 -113 323
rect -79 289 -63 323
rect -129 255 -63 289
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -289 -63 -255
rect -129 -323 -113 -289
rect -79 -323 -63 -289
rect -129 -357 -63 -323
rect -129 -391 -113 -357
rect -79 -391 -63 -357
rect -129 -425 -63 -391
rect -129 -459 -113 -425
rect -79 -459 -63 -425
rect -129 -493 -63 -459
rect -129 -527 -113 -493
rect -79 -527 -63 -493
rect -129 -561 -63 -527
rect -129 -595 -113 -561
rect -79 -595 -63 -561
rect -129 -629 -63 -595
rect -129 -663 -113 -629
rect -79 -663 -63 -629
rect -129 -697 -63 -663
rect -129 -731 -113 -697
rect -79 -731 -63 -697
rect -129 -765 -63 -731
rect -129 -799 -113 -765
rect -79 -799 -63 -765
rect -129 -833 -63 -799
rect -129 -867 -113 -833
rect -79 -867 -63 -833
rect -129 -900 -63 -867
rect -33 867 33 900
rect -33 833 -17 867
rect 17 833 33 867
rect -33 799 33 833
rect -33 765 -17 799
rect 17 765 33 799
rect -33 731 33 765
rect -33 697 -17 731
rect 17 697 33 731
rect -33 663 33 697
rect -33 629 -17 663
rect 17 629 33 663
rect -33 595 33 629
rect -33 561 -17 595
rect 17 561 33 595
rect -33 527 33 561
rect -33 493 -17 527
rect 17 493 33 527
rect -33 459 33 493
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -493 33 -459
rect -33 -527 -17 -493
rect 17 -527 33 -493
rect -33 -561 33 -527
rect -33 -595 -17 -561
rect 17 -595 33 -561
rect -33 -629 33 -595
rect -33 -663 -17 -629
rect 17 -663 33 -629
rect -33 -697 33 -663
rect -33 -731 -17 -697
rect 17 -731 33 -697
rect -33 -765 33 -731
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -833 33 -799
rect -33 -867 -17 -833
rect 17 -867 33 -833
rect -33 -900 33 -867
rect 63 867 129 900
rect 63 833 79 867
rect 113 833 129 867
rect 63 799 129 833
rect 63 765 79 799
rect 113 765 129 799
rect 63 731 129 765
rect 63 697 79 731
rect 113 697 129 731
rect 63 663 129 697
rect 63 629 79 663
rect 113 629 129 663
rect 63 595 129 629
rect 63 561 79 595
rect 113 561 129 595
rect 63 527 129 561
rect 63 493 79 527
rect 113 493 129 527
rect 63 459 129 493
rect 63 425 79 459
rect 113 425 129 459
rect 63 391 129 425
rect 63 357 79 391
rect 113 357 129 391
rect 63 323 129 357
rect 63 289 79 323
rect 113 289 129 323
rect 63 255 129 289
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -289 129 -255
rect 63 -323 79 -289
rect 113 -323 129 -289
rect 63 -357 129 -323
rect 63 -391 79 -357
rect 113 -391 129 -357
rect 63 -425 129 -391
rect 63 -459 79 -425
rect 113 -459 129 -425
rect 63 -493 129 -459
rect 63 -527 79 -493
rect 113 -527 129 -493
rect 63 -561 129 -527
rect 63 -595 79 -561
rect 113 -595 129 -561
rect 63 -629 129 -595
rect 63 -663 79 -629
rect 113 -663 129 -629
rect 63 -697 129 -663
rect 63 -731 79 -697
rect 113 -731 129 -697
rect 63 -765 129 -731
rect 63 -799 79 -765
rect 113 -799 129 -765
rect 63 -833 129 -799
rect 63 -867 79 -833
rect 113 -867 129 -833
rect 63 -900 129 -867
rect 159 867 221 900
rect 159 833 175 867
rect 209 833 221 867
rect 159 799 221 833
rect 159 765 175 799
rect 209 765 221 799
rect 159 731 221 765
rect 159 697 175 731
rect 209 697 221 731
rect 159 663 221 697
rect 159 629 175 663
rect 209 629 221 663
rect 159 595 221 629
rect 159 561 175 595
rect 209 561 221 595
rect 159 527 221 561
rect 159 493 175 527
rect 209 493 221 527
rect 159 459 221 493
rect 159 425 175 459
rect 209 425 221 459
rect 159 391 221 425
rect 159 357 175 391
rect 209 357 221 391
rect 159 323 221 357
rect 159 289 175 323
rect 209 289 221 323
rect 159 255 221 289
rect 159 221 175 255
rect 209 221 221 255
rect 159 187 221 221
rect 159 153 175 187
rect 209 153 221 187
rect 159 119 221 153
rect 159 85 175 119
rect 209 85 221 119
rect 159 51 221 85
rect 159 17 175 51
rect 209 17 221 51
rect 159 -17 221 17
rect 159 -51 175 -17
rect 209 -51 221 -17
rect 159 -85 221 -51
rect 159 -119 175 -85
rect 209 -119 221 -85
rect 159 -153 221 -119
rect 159 -187 175 -153
rect 209 -187 221 -153
rect 159 -221 221 -187
rect 159 -255 175 -221
rect 209 -255 221 -221
rect 159 -289 221 -255
rect 159 -323 175 -289
rect 209 -323 221 -289
rect 159 -357 221 -323
rect 159 -391 175 -357
rect 209 -391 221 -357
rect 159 -425 221 -391
rect 159 -459 175 -425
rect 209 -459 221 -425
rect 159 -493 221 -459
rect 159 -527 175 -493
rect 209 -527 221 -493
rect 159 -561 221 -527
rect 159 -595 175 -561
rect 209 -595 221 -561
rect 159 -629 221 -595
rect 159 -663 175 -629
rect 209 -663 221 -629
rect 159 -697 221 -663
rect 159 -731 175 -697
rect 209 -731 221 -697
rect 159 -765 221 -731
rect 159 -799 175 -765
rect 209 -799 221 -765
rect 159 -833 221 -799
rect 159 -867 175 -833
rect 209 -867 221 -833
rect 159 -900 221 -867
<< pdiffc >>
rect -209 833 -175 867
rect -209 765 -175 799
rect -209 697 -175 731
rect -209 629 -175 663
rect -209 561 -175 595
rect -209 493 -175 527
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -209 -527 -175 -493
rect -209 -595 -175 -561
rect -209 -663 -175 -629
rect -209 -731 -175 -697
rect -209 -799 -175 -765
rect -209 -867 -175 -833
rect -113 833 -79 867
rect -113 765 -79 799
rect -113 697 -79 731
rect -113 629 -79 663
rect -113 561 -79 595
rect -113 493 -79 527
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -113 -527 -79 -493
rect -113 -595 -79 -561
rect -113 -663 -79 -629
rect -113 -731 -79 -697
rect -113 -799 -79 -765
rect -113 -867 -79 -833
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect 79 833 113 867
rect 79 765 113 799
rect 79 697 113 731
rect 79 629 113 663
rect 79 561 113 595
rect 79 493 113 527
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 79 -527 113 -493
rect 79 -595 113 -561
rect 79 -663 113 -629
rect 79 -731 113 -697
rect 79 -799 113 -765
rect 79 -867 113 -833
rect 175 833 209 867
rect 175 765 209 799
rect 175 697 209 731
rect 175 629 209 663
rect 175 561 209 595
rect 175 493 209 527
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
rect 175 -527 209 -493
rect 175 -595 209 -561
rect 175 -663 209 -629
rect 175 -731 209 -697
rect 175 -799 209 -765
rect 175 -867 209 -833
<< nsubdiff >>
rect -323 1049 -221 1083
rect -187 1049 -153 1083
rect -119 1049 -85 1083
rect -51 1049 -17 1083
rect 17 1049 51 1083
rect 85 1049 119 1083
rect 153 1049 187 1083
rect 221 1049 323 1083
rect -323 969 -289 1049
rect -323 901 -289 935
rect 289 969 323 1049
rect 289 901 323 935
rect -323 833 -289 867
rect -323 765 -289 799
rect -323 697 -289 731
rect -323 629 -289 663
rect -323 561 -289 595
rect -323 493 -289 527
rect -323 425 -289 459
rect -323 357 -289 391
rect -323 289 -289 323
rect -323 221 -289 255
rect -323 153 -289 187
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect -323 -187 -289 -153
rect -323 -255 -289 -221
rect -323 -323 -289 -289
rect -323 -391 -289 -357
rect -323 -459 -289 -425
rect -323 -527 -289 -493
rect -323 -595 -289 -561
rect -323 -663 -289 -629
rect -323 -731 -289 -697
rect -323 -799 -289 -765
rect -323 -867 -289 -833
rect 289 833 323 867
rect 289 765 323 799
rect 289 697 323 731
rect 289 629 323 663
rect 289 561 323 595
rect 289 493 323 527
rect 289 425 323 459
rect 289 357 323 391
rect 289 289 323 323
rect 289 221 323 255
rect 289 153 323 187
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect 289 -119 323 -85
rect 289 -187 323 -153
rect 289 -255 323 -221
rect 289 -323 323 -289
rect 289 -391 323 -357
rect 289 -459 323 -425
rect 289 -527 323 -493
rect 289 -595 323 -561
rect 289 -663 323 -629
rect 289 -731 323 -697
rect 289 -799 323 -765
rect 289 -867 323 -833
rect -323 -935 -289 -901
rect -323 -1049 -289 -969
rect 289 -935 323 -901
rect 289 -1049 323 -969
rect -323 -1083 -221 -1049
rect -187 -1083 -153 -1049
rect -119 -1083 -85 -1049
rect -51 -1083 -17 -1049
rect 17 -1083 51 -1049
rect 85 -1083 119 -1049
rect 153 -1083 187 -1049
rect 221 -1083 323 -1049
<< nsubdiffcont >>
rect -221 1049 -187 1083
rect -153 1049 -119 1083
rect -85 1049 -51 1083
rect -17 1049 17 1083
rect 51 1049 85 1083
rect 119 1049 153 1083
rect 187 1049 221 1083
rect -323 935 -289 969
rect 289 935 323 969
rect -323 867 -289 901
rect -323 799 -289 833
rect -323 731 -289 765
rect -323 663 -289 697
rect -323 595 -289 629
rect -323 527 -289 561
rect -323 459 -289 493
rect -323 391 -289 425
rect -323 323 -289 357
rect -323 255 -289 289
rect -323 187 -289 221
rect -323 119 -289 153
rect -323 51 -289 85
rect -323 -17 -289 17
rect -323 -85 -289 -51
rect -323 -153 -289 -119
rect -323 -221 -289 -187
rect -323 -289 -289 -255
rect -323 -357 -289 -323
rect -323 -425 -289 -391
rect -323 -493 -289 -459
rect -323 -561 -289 -527
rect -323 -629 -289 -595
rect -323 -697 -289 -663
rect -323 -765 -289 -731
rect -323 -833 -289 -799
rect -323 -901 -289 -867
rect 289 867 323 901
rect 289 799 323 833
rect 289 731 323 765
rect 289 663 323 697
rect 289 595 323 629
rect 289 527 323 561
rect 289 459 323 493
rect 289 391 323 425
rect 289 323 323 357
rect 289 255 323 289
rect 289 187 323 221
rect 289 119 323 153
rect 289 51 323 85
rect 289 -17 323 17
rect 289 -85 323 -51
rect 289 -153 323 -119
rect 289 -221 323 -187
rect 289 -289 323 -255
rect 289 -357 323 -323
rect 289 -425 323 -391
rect 289 -493 323 -459
rect 289 -561 323 -527
rect 289 -629 323 -595
rect 289 -697 323 -663
rect 289 -765 323 -731
rect 289 -833 323 -799
rect 289 -901 323 -867
rect -323 -969 -289 -935
rect 289 -969 323 -935
rect -221 -1083 -187 -1049
rect -153 -1083 -119 -1049
rect -85 -1083 -51 -1049
rect -17 -1083 17 -1049
rect 51 -1083 85 -1049
rect 119 -1083 153 -1049
rect 187 -1083 221 -1049
<< poly >>
rect -81 981 -15 997
rect -81 947 -65 981
rect -31 947 -15 981
rect -81 931 -15 947
rect 111 981 177 997
rect 111 947 127 981
rect 161 947 177 981
rect 111 931 177 947
rect -159 900 -129 926
rect -63 900 -33 931
rect 33 900 63 926
rect 129 900 159 931
rect -159 -931 -129 -900
rect -63 -926 -33 -900
rect 33 -931 63 -900
rect 129 -926 159 -900
rect -177 -947 -111 -931
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect -177 -997 -111 -981
rect 15 -947 81 -931
rect 15 -981 31 -947
rect 65 -981 81 -947
rect 15 -997 81 -981
<< polycont >>
rect -65 947 -31 981
rect 127 947 161 981
rect -161 -981 -127 -947
rect 31 -981 65 -947
<< locali >>
rect -323 1049 -221 1083
rect -187 1049 -153 1083
rect -119 1049 -85 1083
rect -51 1049 -17 1083
rect 17 1049 51 1083
rect 85 1049 119 1083
rect 153 1049 187 1083
rect 221 1049 323 1083
rect -323 969 -289 1049
rect -81 947 -65 981
rect -31 947 -15 981
rect 111 947 127 981
rect 161 947 177 981
rect 289 969 323 1049
rect -323 901 -289 935
rect -323 833 -289 867
rect -323 765 -289 799
rect -323 697 -289 731
rect -323 629 -289 663
rect -323 561 -289 595
rect -323 493 -289 527
rect -323 425 -289 459
rect -323 357 -289 391
rect -323 289 -289 323
rect -323 221 -289 255
rect -323 153 -289 187
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect -323 -187 -289 -153
rect -323 -255 -289 -221
rect -323 -323 -289 -289
rect -323 -391 -289 -357
rect -323 -459 -289 -425
rect -323 -527 -289 -493
rect -323 -595 -289 -561
rect -323 -663 -289 -629
rect -323 -731 -289 -697
rect -323 -799 -289 -765
rect -323 -867 -289 -833
rect -323 -935 -289 -901
rect -209 881 -175 904
rect -209 809 -175 833
rect -209 737 -175 765
rect -209 665 -175 697
rect -209 595 -175 629
rect -209 527 -175 559
rect -209 459 -175 487
rect -209 391 -175 415
rect -209 323 -175 343
rect -209 255 -175 271
rect -209 187 -175 199
rect -209 119 -175 127
rect -209 51 -175 55
rect -209 -55 -175 -51
rect -209 -127 -175 -119
rect -209 -199 -175 -187
rect -209 -271 -175 -255
rect -209 -343 -175 -323
rect -209 -415 -175 -391
rect -209 -487 -175 -459
rect -209 -559 -175 -527
rect -209 -629 -175 -595
rect -209 -697 -175 -665
rect -209 -765 -175 -737
rect -209 -833 -175 -809
rect -209 -904 -175 -881
rect -113 881 -79 904
rect -113 809 -79 833
rect -113 737 -79 765
rect -113 665 -79 697
rect -113 595 -79 629
rect -113 527 -79 559
rect -113 459 -79 487
rect -113 391 -79 415
rect -113 323 -79 343
rect -113 255 -79 271
rect -113 187 -79 199
rect -113 119 -79 127
rect -113 51 -79 55
rect -113 -55 -79 -51
rect -113 -127 -79 -119
rect -113 -199 -79 -187
rect -113 -271 -79 -255
rect -113 -343 -79 -323
rect -113 -415 -79 -391
rect -113 -487 -79 -459
rect -113 -559 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -665
rect -113 -765 -79 -737
rect -113 -833 -79 -809
rect -113 -904 -79 -881
rect -17 881 17 904
rect -17 809 17 833
rect -17 737 17 765
rect -17 665 17 697
rect -17 595 17 629
rect -17 527 17 559
rect -17 459 17 487
rect -17 391 17 415
rect -17 323 17 343
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -343 17 -323
rect -17 -415 17 -391
rect -17 -487 17 -459
rect -17 -559 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -665
rect -17 -765 17 -737
rect -17 -833 17 -809
rect -17 -904 17 -881
rect 79 881 113 904
rect 79 809 113 833
rect 79 737 113 765
rect 79 665 113 697
rect 79 595 113 629
rect 79 527 113 559
rect 79 459 113 487
rect 79 391 113 415
rect 79 323 113 343
rect 79 255 113 271
rect 79 187 113 199
rect 79 119 113 127
rect 79 51 113 55
rect 79 -55 113 -51
rect 79 -127 113 -119
rect 79 -199 113 -187
rect 79 -271 113 -255
rect 79 -343 113 -323
rect 79 -415 113 -391
rect 79 -487 113 -459
rect 79 -559 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -665
rect 79 -765 113 -737
rect 79 -833 113 -809
rect 79 -904 113 -881
rect 175 881 209 904
rect 175 809 209 833
rect 175 737 209 765
rect 175 665 209 697
rect 175 595 209 629
rect 175 527 209 559
rect 175 459 209 487
rect 175 391 209 415
rect 175 323 209 343
rect 175 255 209 271
rect 175 187 209 199
rect 175 119 209 127
rect 175 51 209 55
rect 175 -55 209 -51
rect 175 -127 209 -119
rect 175 -199 209 -187
rect 175 -271 209 -255
rect 175 -343 209 -323
rect 175 -415 209 -391
rect 175 -487 209 -459
rect 175 -559 209 -527
rect 175 -629 209 -595
rect 175 -697 209 -665
rect 175 -765 209 -737
rect 175 -833 209 -809
rect 175 -904 209 -881
rect 289 901 323 935
rect 289 833 323 867
rect 289 765 323 799
rect 289 697 323 731
rect 289 629 323 663
rect 289 561 323 595
rect 289 493 323 527
rect 289 425 323 459
rect 289 357 323 391
rect 289 289 323 323
rect 289 221 323 255
rect 289 153 323 187
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect 289 -119 323 -85
rect 289 -187 323 -153
rect 289 -255 323 -221
rect 289 -323 323 -289
rect 289 -391 323 -357
rect 289 -459 323 -425
rect 289 -527 323 -493
rect 289 -595 323 -561
rect 289 -663 323 -629
rect 289 -731 323 -697
rect 289 -799 323 -765
rect 289 -867 323 -833
rect 289 -935 323 -901
rect -323 -1049 -289 -969
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect 15 -981 31 -947
rect 65 -981 81 -947
rect 289 -1049 323 -969
rect -323 -1083 -221 -1049
rect -187 -1083 -153 -1049
rect -119 -1083 -85 -1049
rect -51 -1083 -17 -1049
rect 17 -1083 51 -1049
rect 85 -1083 119 -1049
rect 153 -1083 187 -1049
rect 221 -1083 323 -1049
<< viali >>
rect -65 947 -31 981
rect 127 947 161 981
rect -209 867 -175 881
rect -209 847 -175 867
rect -209 799 -175 809
rect -209 775 -175 799
rect -209 731 -175 737
rect -209 703 -175 731
rect -209 663 -175 665
rect -209 631 -175 663
rect -209 561 -175 593
rect -209 559 -175 561
rect -209 493 -175 521
rect -209 487 -175 493
rect -209 425 -175 449
rect -209 415 -175 425
rect -209 357 -175 377
rect -209 343 -175 357
rect -209 289 -175 305
rect -209 271 -175 289
rect -209 221 -175 233
rect -209 199 -175 221
rect -209 153 -175 161
rect -209 127 -175 153
rect -209 85 -175 89
rect -209 55 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -55
rect -209 -89 -175 -85
rect -209 -153 -175 -127
rect -209 -161 -175 -153
rect -209 -221 -175 -199
rect -209 -233 -175 -221
rect -209 -289 -175 -271
rect -209 -305 -175 -289
rect -209 -357 -175 -343
rect -209 -377 -175 -357
rect -209 -425 -175 -415
rect -209 -449 -175 -425
rect -209 -493 -175 -487
rect -209 -521 -175 -493
rect -209 -561 -175 -559
rect -209 -593 -175 -561
rect -209 -663 -175 -631
rect -209 -665 -175 -663
rect -209 -731 -175 -703
rect -209 -737 -175 -731
rect -209 -799 -175 -775
rect -209 -809 -175 -799
rect -209 -867 -175 -847
rect -209 -881 -175 -867
rect -113 867 -79 881
rect -113 847 -79 867
rect -113 799 -79 809
rect -113 775 -79 799
rect -113 731 -79 737
rect -113 703 -79 731
rect -113 663 -79 665
rect -113 631 -79 663
rect -113 561 -79 593
rect -113 559 -79 561
rect -113 493 -79 521
rect -113 487 -79 493
rect -113 425 -79 449
rect -113 415 -79 425
rect -113 357 -79 377
rect -113 343 -79 357
rect -113 289 -79 305
rect -113 271 -79 289
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -113 -289 -79 -271
rect -113 -305 -79 -289
rect -113 -357 -79 -343
rect -113 -377 -79 -357
rect -113 -425 -79 -415
rect -113 -449 -79 -425
rect -113 -493 -79 -487
rect -113 -521 -79 -493
rect -113 -561 -79 -559
rect -113 -593 -79 -561
rect -113 -663 -79 -631
rect -113 -665 -79 -663
rect -113 -731 -79 -703
rect -113 -737 -79 -731
rect -113 -799 -79 -775
rect -113 -809 -79 -799
rect -113 -867 -79 -847
rect -113 -881 -79 -867
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect 79 867 113 881
rect 79 847 113 867
rect 79 799 113 809
rect 79 775 113 799
rect 79 731 113 737
rect 79 703 113 731
rect 79 663 113 665
rect 79 631 113 663
rect 79 561 113 593
rect 79 559 113 561
rect 79 493 113 521
rect 79 487 113 493
rect 79 425 113 449
rect 79 415 113 425
rect 79 357 113 377
rect 79 343 113 357
rect 79 289 113 305
rect 79 271 113 289
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
rect 79 -289 113 -271
rect 79 -305 113 -289
rect 79 -357 113 -343
rect 79 -377 113 -357
rect 79 -425 113 -415
rect 79 -449 113 -425
rect 79 -493 113 -487
rect 79 -521 113 -493
rect 79 -561 113 -559
rect 79 -593 113 -561
rect 79 -663 113 -631
rect 79 -665 113 -663
rect 79 -731 113 -703
rect 79 -737 113 -731
rect 79 -799 113 -775
rect 79 -809 113 -799
rect 79 -867 113 -847
rect 79 -881 113 -867
rect 175 867 209 881
rect 175 847 209 867
rect 175 799 209 809
rect 175 775 209 799
rect 175 731 209 737
rect 175 703 209 731
rect 175 663 209 665
rect 175 631 209 663
rect 175 561 209 593
rect 175 559 209 561
rect 175 493 209 521
rect 175 487 209 493
rect 175 425 209 449
rect 175 415 209 425
rect 175 357 209 377
rect 175 343 209 357
rect 175 289 209 305
rect 175 271 209 289
rect 175 221 209 233
rect 175 199 209 221
rect 175 153 209 161
rect 175 127 209 153
rect 175 85 209 89
rect 175 55 209 85
rect 175 -17 209 17
rect 175 -85 209 -55
rect 175 -89 209 -85
rect 175 -153 209 -127
rect 175 -161 209 -153
rect 175 -221 209 -199
rect 175 -233 209 -221
rect 175 -289 209 -271
rect 175 -305 209 -289
rect 175 -357 209 -343
rect 175 -377 209 -357
rect 175 -425 209 -415
rect 175 -449 209 -425
rect 175 -493 209 -487
rect 175 -521 209 -493
rect 175 -561 209 -559
rect 175 -593 209 -561
rect 175 -663 209 -631
rect 175 -665 209 -663
rect 175 -731 209 -703
rect 175 -737 209 -731
rect 175 -799 209 -775
rect 175 -809 209 -799
rect 175 -867 209 -847
rect 175 -881 209 -867
rect -161 -981 -127 -947
rect 31 -981 65 -947
<< metal1 >>
rect -77 981 -19 987
rect -77 947 -65 981
rect -31 947 -19 981
rect -77 941 -19 947
rect 115 981 173 987
rect 115 947 127 981
rect 161 947 173 981
rect 115 941 173 947
rect -215 881 -169 900
rect -215 847 -209 881
rect -175 847 -169 881
rect -215 809 -169 847
rect -215 775 -209 809
rect -175 775 -169 809
rect -215 737 -169 775
rect -215 703 -209 737
rect -175 703 -169 737
rect -215 665 -169 703
rect -215 631 -209 665
rect -175 631 -169 665
rect -215 593 -169 631
rect -215 559 -209 593
rect -175 559 -169 593
rect -215 521 -169 559
rect -215 487 -209 521
rect -175 487 -169 521
rect -215 449 -169 487
rect -215 415 -209 449
rect -175 415 -169 449
rect -215 377 -169 415
rect -215 343 -209 377
rect -175 343 -169 377
rect -215 305 -169 343
rect -215 271 -209 305
rect -175 271 -169 305
rect -215 233 -169 271
rect -215 199 -209 233
rect -175 199 -169 233
rect -215 161 -169 199
rect -215 127 -209 161
rect -175 127 -169 161
rect -215 89 -169 127
rect -215 55 -209 89
rect -175 55 -169 89
rect -215 17 -169 55
rect -215 -17 -209 17
rect -175 -17 -169 17
rect -215 -55 -169 -17
rect -215 -89 -209 -55
rect -175 -89 -169 -55
rect -215 -127 -169 -89
rect -215 -161 -209 -127
rect -175 -161 -169 -127
rect -215 -199 -169 -161
rect -215 -233 -209 -199
rect -175 -233 -169 -199
rect -215 -271 -169 -233
rect -215 -305 -209 -271
rect -175 -305 -169 -271
rect -215 -343 -169 -305
rect -215 -377 -209 -343
rect -175 -377 -169 -343
rect -215 -415 -169 -377
rect -215 -449 -209 -415
rect -175 -449 -169 -415
rect -215 -487 -169 -449
rect -215 -521 -209 -487
rect -175 -521 -169 -487
rect -215 -559 -169 -521
rect -215 -593 -209 -559
rect -175 -593 -169 -559
rect -215 -631 -169 -593
rect -215 -665 -209 -631
rect -175 -665 -169 -631
rect -215 -703 -169 -665
rect -215 -737 -209 -703
rect -175 -737 -169 -703
rect -215 -775 -169 -737
rect -215 -809 -209 -775
rect -175 -809 -169 -775
rect -215 -847 -169 -809
rect -215 -881 -209 -847
rect -175 -881 -169 -847
rect -215 -900 -169 -881
rect -119 881 -73 900
rect -119 847 -113 881
rect -79 847 -73 881
rect -119 809 -73 847
rect -119 775 -113 809
rect -79 775 -73 809
rect -119 737 -73 775
rect -119 703 -113 737
rect -79 703 -73 737
rect -119 665 -73 703
rect -119 631 -113 665
rect -79 631 -73 665
rect -119 593 -73 631
rect -119 559 -113 593
rect -79 559 -73 593
rect -119 521 -73 559
rect -119 487 -113 521
rect -79 487 -73 521
rect -119 449 -73 487
rect -119 415 -113 449
rect -79 415 -73 449
rect -119 377 -73 415
rect -119 343 -113 377
rect -79 343 -73 377
rect -119 305 -73 343
rect -119 271 -113 305
rect -79 271 -73 305
rect -119 233 -73 271
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -271 -73 -233
rect -119 -305 -113 -271
rect -79 -305 -73 -271
rect -119 -343 -73 -305
rect -119 -377 -113 -343
rect -79 -377 -73 -343
rect -119 -415 -73 -377
rect -119 -449 -113 -415
rect -79 -449 -73 -415
rect -119 -487 -73 -449
rect -119 -521 -113 -487
rect -79 -521 -73 -487
rect -119 -559 -73 -521
rect -119 -593 -113 -559
rect -79 -593 -73 -559
rect -119 -631 -73 -593
rect -119 -665 -113 -631
rect -79 -665 -73 -631
rect -119 -703 -73 -665
rect -119 -737 -113 -703
rect -79 -737 -73 -703
rect -119 -775 -73 -737
rect -119 -809 -113 -775
rect -79 -809 -73 -775
rect -119 -847 -73 -809
rect -119 -881 -113 -847
rect -79 -881 -73 -847
rect -119 -900 -73 -881
rect -23 881 23 900
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -900 23 -881
rect 73 881 119 900
rect 73 847 79 881
rect 113 847 119 881
rect 73 809 119 847
rect 73 775 79 809
rect 113 775 119 809
rect 73 737 119 775
rect 73 703 79 737
rect 113 703 119 737
rect 73 665 119 703
rect 73 631 79 665
rect 113 631 119 665
rect 73 593 119 631
rect 73 559 79 593
rect 113 559 119 593
rect 73 521 119 559
rect 73 487 79 521
rect 113 487 119 521
rect 73 449 119 487
rect 73 415 79 449
rect 113 415 119 449
rect 73 377 119 415
rect 73 343 79 377
rect 113 343 119 377
rect 73 305 119 343
rect 73 271 79 305
rect 113 271 119 305
rect 73 233 119 271
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -271 119 -233
rect 73 -305 79 -271
rect 113 -305 119 -271
rect 73 -343 119 -305
rect 73 -377 79 -343
rect 113 -377 119 -343
rect 73 -415 119 -377
rect 73 -449 79 -415
rect 113 -449 119 -415
rect 73 -487 119 -449
rect 73 -521 79 -487
rect 113 -521 119 -487
rect 73 -559 119 -521
rect 73 -593 79 -559
rect 113 -593 119 -559
rect 73 -631 119 -593
rect 73 -665 79 -631
rect 113 -665 119 -631
rect 73 -703 119 -665
rect 73 -737 79 -703
rect 113 -737 119 -703
rect 73 -775 119 -737
rect 73 -809 79 -775
rect 113 -809 119 -775
rect 73 -847 119 -809
rect 73 -881 79 -847
rect 113 -881 119 -847
rect 73 -900 119 -881
rect 169 881 215 900
rect 169 847 175 881
rect 209 847 215 881
rect 169 809 215 847
rect 169 775 175 809
rect 209 775 215 809
rect 169 737 215 775
rect 169 703 175 737
rect 209 703 215 737
rect 169 665 215 703
rect 169 631 175 665
rect 209 631 215 665
rect 169 593 215 631
rect 169 559 175 593
rect 209 559 215 593
rect 169 521 215 559
rect 169 487 175 521
rect 209 487 215 521
rect 169 449 215 487
rect 169 415 175 449
rect 209 415 215 449
rect 169 377 215 415
rect 169 343 175 377
rect 209 343 215 377
rect 169 305 215 343
rect 169 271 175 305
rect 209 271 215 305
rect 169 233 215 271
rect 169 199 175 233
rect 209 199 215 233
rect 169 161 215 199
rect 169 127 175 161
rect 209 127 215 161
rect 169 89 215 127
rect 169 55 175 89
rect 209 55 215 89
rect 169 17 215 55
rect 169 -17 175 17
rect 209 -17 215 17
rect 169 -55 215 -17
rect 169 -89 175 -55
rect 209 -89 215 -55
rect 169 -127 215 -89
rect 169 -161 175 -127
rect 209 -161 215 -127
rect 169 -199 215 -161
rect 169 -233 175 -199
rect 209 -233 215 -199
rect 169 -271 215 -233
rect 169 -305 175 -271
rect 209 -305 215 -271
rect 169 -343 215 -305
rect 169 -377 175 -343
rect 209 -377 215 -343
rect 169 -415 215 -377
rect 169 -449 175 -415
rect 209 -449 215 -415
rect 169 -487 215 -449
rect 169 -521 175 -487
rect 209 -521 215 -487
rect 169 -559 215 -521
rect 169 -593 175 -559
rect 209 -593 215 -559
rect 169 -631 215 -593
rect 169 -665 175 -631
rect 209 -665 215 -631
rect 169 -703 215 -665
rect 169 -737 175 -703
rect 209 -737 215 -703
rect 169 -775 215 -737
rect 169 -809 175 -775
rect 209 -809 215 -775
rect 169 -847 215 -809
rect 169 -881 175 -847
rect 209 -881 215 -847
rect 169 -900 215 -881
rect -173 -947 -115 -941
rect -173 -981 -161 -947
rect -127 -981 -115 -947
rect -173 -987 -115 -981
rect 19 -947 77 -941
rect 19 -981 31 -947
rect 65 -981 77 -947
rect 19 -987 77 -981
<< properties >>
string FIXED_BBOX -306 -1066 306 1066
<< end >>
