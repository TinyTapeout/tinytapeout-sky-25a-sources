magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 832 240
<< ntap >>
rect -48 60 880 100
rect -48 100 880 140
rect -48 140 880 180
rect -48 180 48 220
rect 784 180 880 220
rect -48 220 48 260
rect 784 220 880 260
<< locali >>
rect -48 60 880 100
rect -48 100 880 140
rect -48 140 880 180
rect -48 180 48 220
rect 784 180 880 220
rect -48 220 48 260
rect 784 220 880 260
<< ntapc >>
rect 80 100 720 140
<< nwell >>
rect -92 -64 924 304
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 832 240
<< end >>
