magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -78 1981 -20 1987
rect 118 1981 176 1987
rect -78 1947 -66 1981
rect 118 1947 130 1981
rect -78 1941 -20 1947
rect 118 1941 176 1947
rect -176 -1947 -118 -1941
rect 20 -1947 78 -1941
rect -176 -1981 -164 -1947
rect 20 -1981 32 -1947
rect -176 -1987 -118 -1981
rect 20 -1987 78 -1981
<< nwell >>
rect -363 -2119 363 2119
<< pmos >>
rect -167 -1900 -127 1900
rect -69 -1900 -29 1900
rect 29 -1900 69 1900
rect 127 -1900 167 1900
<< pdiff >>
rect -225 1887 -167 1900
rect -225 1853 -213 1887
rect -179 1853 -167 1887
rect -225 1819 -167 1853
rect -225 1785 -213 1819
rect -179 1785 -167 1819
rect -225 1751 -167 1785
rect -225 1717 -213 1751
rect -179 1717 -167 1751
rect -225 1683 -167 1717
rect -225 1649 -213 1683
rect -179 1649 -167 1683
rect -225 1615 -167 1649
rect -225 1581 -213 1615
rect -179 1581 -167 1615
rect -225 1547 -167 1581
rect -225 1513 -213 1547
rect -179 1513 -167 1547
rect -225 1479 -167 1513
rect -225 1445 -213 1479
rect -179 1445 -167 1479
rect -225 1411 -167 1445
rect -225 1377 -213 1411
rect -179 1377 -167 1411
rect -225 1343 -167 1377
rect -225 1309 -213 1343
rect -179 1309 -167 1343
rect -225 1275 -167 1309
rect -225 1241 -213 1275
rect -179 1241 -167 1275
rect -225 1207 -167 1241
rect -225 1173 -213 1207
rect -179 1173 -167 1207
rect -225 1139 -167 1173
rect -225 1105 -213 1139
rect -179 1105 -167 1139
rect -225 1071 -167 1105
rect -225 1037 -213 1071
rect -179 1037 -167 1071
rect -225 1003 -167 1037
rect -225 969 -213 1003
rect -179 969 -167 1003
rect -225 935 -167 969
rect -225 901 -213 935
rect -179 901 -167 935
rect -225 867 -167 901
rect -225 833 -213 867
rect -179 833 -167 867
rect -225 799 -167 833
rect -225 765 -213 799
rect -179 765 -167 799
rect -225 731 -167 765
rect -225 697 -213 731
rect -179 697 -167 731
rect -225 663 -167 697
rect -225 629 -213 663
rect -179 629 -167 663
rect -225 595 -167 629
rect -225 561 -213 595
rect -179 561 -167 595
rect -225 527 -167 561
rect -225 493 -213 527
rect -179 493 -167 527
rect -225 459 -167 493
rect -225 425 -213 459
rect -179 425 -167 459
rect -225 391 -167 425
rect -225 357 -213 391
rect -179 357 -167 391
rect -225 323 -167 357
rect -225 289 -213 323
rect -179 289 -167 323
rect -225 255 -167 289
rect -225 221 -213 255
rect -179 221 -167 255
rect -225 187 -167 221
rect -225 153 -213 187
rect -179 153 -167 187
rect -225 119 -167 153
rect -225 85 -213 119
rect -179 85 -167 119
rect -225 51 -167 85
rect -225 17 -213 51
rect -179 17 -167 51
rect -225 -17 -167 17
rect -225 -51 -213 -17
rect -179 -51 -167 -17
rect -225 -85 -167 -51
rect -225 -119 -213 -85
rect -179 -119 -167 -85
rect -225 -153 -167 -119
rect -225 -187 -213 -153
rect -179 -187 -167 -153
rect -225 -221 -167 -187
rect -225 -255 -213 -221
rect -179 -255 -167 -221
rect -225 -289 -167 -255
rect -225 -323 -213 -289
rect -179 -323 -167 -289
rect -225 -357 -167 -323
rect -225 -391 -213 -357
rect -179 -391 -167 -357
rect -225 -425 -167 -391
rect -225 -459 -213 -425
rect -179 -459 -167 -425
rect -225 -493 -167 -459
rect -225 -527 -213 -493
rect -179 -527 -167 -493
rect -225 -561 -167 -527
rect -225 -595 -213 -561
rect -179 -595 -167 -561
rect -225 -629 -167 -595
rect -225 -663 -213 -629
rect -179 -663 -167 -629
rect -225 -697 -167 -663
rect -225 -731 -213 -697
rect -179 -731 -167 -697
rect -225 -765 -167 -731
rect -225 -799 -213 -765
rect -179 -799 -167 -765
rect -225 -833 -167 -799
rect -225 -867 -213 -833
rect -179 -867 -167 -833
rect -225 -901 -167 -867
rect -225 -935 -213 -901
rect -179 -935 -167 -901
rect -225 -969 -167 -935
rect -225 -1003 -213 -969
rect -179 -1003 -167 -969
rect -225 -1037 -167 -1003
rect -225 -1071 -213 -1037
rect -179 -1071 -167 -1037
rect -225 -1105 -167 -1071
rect -225 -1139 -213 -1105
rect -179 -1139 -167 -1105
rect -225 -1173 -167 -1139
rect -225 -1207 -213 -1173
rect -179 -1207 -167 -1173
rect -225 -1241 -167 -1207
rect -225 -1275 -213 -1241
rect -179 -1275 -167 -1241
rect -225 -1309 -167 -1275
rect -225 -1343 -213 -1309
rect -179 -1343 -167 -1309
rect -225 -1377 -167 -1343
rect -225 -1411 -213 -1377
rect -179 -1411 -167 -1377
rect -225 -1445 -167 -1411
rect -225 -1479 -213 -1445
rect -179 -1479 -167 -1445
rect -225 -1513 -167 -1479
rect -225 -1547 -213 -1513
rect -179 -1547 -167 -1513
rect -225 -1581 -167 -1547
rect -225 -1615 -213 -1581
rect -179 -1615 -167 -1581
rect -225 -1649 -167 -1615
rect -225 -1683 -213 -1649
rect -179 -1683 -167 -1649
rect -225 -1717 -167 -1683
rect -225 -1751 -213 -1717
rect -179 -1751 -167 -1717
rect -225 -1785 -167 -1751
rect -225 -1819 -213 -1785
rect -179 -1819 -167 -1785
rect -225 -1853 -167 -1819
rect -225 -1887 -213 -1853
rect -179 -1887 -167 -1853
rect -225 -1900 -167 -1887
rect -127 1887 -69 1900
rect -127 1853 -115 1887
rect -81 1853 -69 1887
rect -127 1819 -69 1853
rect -127 1785 -115 1819
rect -81 1785 -69 1819
rect -127 1751 -69 1785
rect -127 1717 -115 1751
rect -81 1717 -69 1751
rect -127 1683 -69 1717
rect -127 1649 -115 1683
rect -81 1649 -69 1683
rect -127 1615 -69 1649
rect -127 1581 -115 1615
rect -81 1581 -69 1615
rect -127 1547 -69 1581
rect -127 1513 -115 1547
rect -81 1513 -69 1547
rect -127 1479 -69 1513
rect -127 1445 -115 1479
rect -81 1445 -69 1479
rect -127 1411 -69 1445
rect -127 1377 -115 1411
rect -81 1377 -69 1411
rect -127 1343 -69 1377
rect -127 1309 -115 1343
rect -81 1309 -69 1343
rect -127 1275 -69 1309
rect -127 1241 -115 1275
rect -81 1241 -69 1275
rect -127 1207 -69 1241
rect -127 1173 -115 1207
rect -81 1173 -69 1207
rect -127 1139 -69 1173
rect -127 1105 -115 1139
rect -81 1105 -69 1139
rect -127 1071 -69 1105
rect -127 1037 -115 1071
rect -81 1037 -69 1071
rect -127 1003 -69 1037
rect -127 969 -115 1003
rect -81 969 -69 1003
rect -127 935 -69 969
rect -127 901 -115 935
rect -81 901 -69 935
rect -127 867 -69 901
rect -127 833 -115 867
rect -81 833 -69 867
rect -127 799 -69 833
rect -127 765 -115 799
rect -81 765 -69 799
rect -127 731 -69 765
rect -127 697 -115 731
rect -81 697 -69 731
rect -127 663 -69 697
rect -127 629 -115 663
rect -81 629 -69 663
rect -127 595 -69 629
rect -127 561 -115 595
rect -81 561 -69 595
rect -127 527 -69 561
rect -127 493 -115 527
rect -81 493 -69 527
rect -127 459 -69 493
rect -127 425 -115 459
rect -81 425 -69 459
rect -127 391 -69 425
rect -127 357 -115 391
rect -81 357 -69 391
rect -127 323 -69 357
rect -127 289 -115 323
rect -81 289 -69 323
rect -127 255 -69 289
rect -127 221 -115 255
rect -81 221 -69 255
rect -127 187 -69 221
rect -127 153 -115 187
rect -81 153 -69 187
rect -127 119 -69 153
rect -127 85 -115 119
rect -81 85 -69 119
rect -127 51 -69 85
rect -127 17 -115 51
rect -81 17 -69 51
rect -127 -17 -69 17
rect -127 -51 -115 -17
rect -81 -51 -69 -17
rect -127 -85 -69 -51
rect -127 -119 -115 -85
rect -81 -119 -69 -85
rect -127 -153 -69 -119
rect -127 -187 -115 -153
rect -81 -187 -69 -153
rect -127 -221 -69 -187
rect -127 -255 -115 -221
rect -81 -255 -69 -221
rect -127 -289 -69 -255
rect -127 -323 -115 -289
rect -81 -323 -69 -289
rect -127 -357 -69 -323
rect -127 -391 -115 -357
rect -81 -391 -69 -357
rect -127 -425 -69 -391
rect -127 -459 -115 -425
rect -81 -459 -69 -425
rect -127 -493 -69 -459
rect -127 -527 -115 -493
rect -81 -527 -69 -493
rect -127 -561 -69 -527
rect -127 -595 -115 -561
rect -81 -595 -69 -561
rect -127 -629 -69 -595
rect -127 -663 -115 -629
rect -81 -663 -69 -629
rect -127 -697 -69 -663
rect -127 -731 -115 -697
rect -81 -731 -69 -697
rect -127 -765 -69 -731
rect -127 -799 -115 -765
rect -81 -799 -69 -765
rect -127 -833 -69 -799
rect -127 -867 -115 -833
rect -81 -867 -69 -833
rect -127 -901 -69 -867
rect -127 -935 -115 -901
rect -81 -935 -69 -901
rect -127 -969 -69 -935
rect -127 -1003 -115 -969
rect -81 -1003 -69 -969
rect -127 -1037 -69 -1003
rect -127 -1071 -115 -1037
rect -81 -1071 -69 -1037
rect -127 -1105 -69 -1071
rect -127 -1139 -115 -1105
rect -81 -1139 -69 -1105
rect -127 -1173 -69 -1139
rect -127 -1207 -115 -1173
rect -81 -1207 -69 -1173
rect -127 -1241 -69 -1207
rect -127 -1275 -115 -1241
rect -81 -1275 -69 -1241
rect -127 -1309 -69 -1275
rect -127 -1343 -115 -1309
rect -81 -1343 -69 -1309
rect -127 -1377 -69 -1343
rect -127 -1411 -115 -1377
rect -81 -1411 -69 -1377
rect -127 -1445 -69 -1411
rect -127 -1479 -115 -1445
rect -81 -1479 -69 -1445
rect -127 -1513 -69 -1479
rect -127 -1547 -115 -1513
rect -81 -1547 -69 -1513
rect -127 -1581 -69 -1547
rect -127 -1615 -115 -1581
rect -81 -1615 -69 -1581
rect -127 -1649 -69 -1615
rect -127 -1683 -115 -1649
rect -81 -1683 -69 -1649
rect -127 -1717 -69 -1683
rect -127 -1751 -115 -1717
rect -81 -1751 -69 -1717
rect -127 -1785 -69 -1751
rect -127 -1819 -115 -1785
rect -81 -1819 -69 -1785
rect -127 -1853 -69 -1819
rect -127 -1887 -115 -1853
rect -81 -1887 -69 -1853
rect -127 -1900 -69 -1887
rect -29 1887 29 1900
rect -29 1853 -17 1887
rect 17 1853 29 1887
rect -29 1819 29 1853
rect -29 1785 -17 1819
rect 17 1785 29 1819
rect -29 1751 29 1785
rect -29 1717 -17 1751
rect 17 1717 29 1751
rect -29 1683 29 1717
rect -29 1649 -17 1683
rect 17 1649 29 1683
rect -29 1615 29 1649
rect -29 1581 -17 1615
rect 17 1581 29 1615
rect -29 1547 29 1581
rect -29 1513 -17 1547
rect 17 1513 29 1547
rect -29 1479 29 1513
rect -29 1445 -17 1479
rect 17 1445 29 1479
rect -29 1411 29 1445
rect -29 1377 -17 1411
rect 17 1377 29 1411
rect -29 1343 29 1377
rect -29 1309 -17 1343
rect 17 1309 29 1343
rect -29 1275 29 1309
rect -29 1241 -17 1275
rect 17 1241 29 1275
rect -29 1207 29 1241
rect -29 1173 -17 1207
rect 17 1173 29 1207
rect -29 1139 29 1173
rect -29 1105 -17 1139
rect 17 1105 29 1139
rect -29 1071 29 1105
rect -29 1037 -17 1071
rect 17 1037 29 1071
rect -29 1003 29 1037
rect -29 969 -17 1003
rect 17 969 29 1003
rect -29 935 29 969
rect -29 901 -17 935
rect 17 901 29 935
rect -29 867 29 901
rect -29 833 -17 867
rect 17 833 29 867
rect -29 799 29 833
rect -29 765 -17 799
rect 17 765 29 799
rect -29 731 29 765
rect -29 697 -17 731
rect 17 697 29 731
rect -29 663 29 697
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -697 29 -663
rect -29 -731 -17 -697
rect 17 -731 29 -697
rect -29 -765 29 -731
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -833 29 -799
rect -29 -867 -17 -833
rect 17 -867 29 -833
rect -29 -901 29 -867
rect -29 -935 -17 -901
rect 17 -935 29 -901
rect -29 -969 29 -935
rect -29 -1003 -17 -969
rect 17 -1003 29 -969
rect -29 -1037 29 -1003
rect -29 -1071 -17 -1037
rect 17 -1071 29 -1037
rect -29 -1105 29 -1071
rect -29 -1139 -17 -1105
rect 17 -1139 29 -1105
rect -29 -1173 29 -1139
rect -29 -1207 -17 -1173
rect 17 -1207 29 -1173
rect -29 -1241 29 -1207
rect -29 -1275 -17 -1241
rect 17 -1275 29 -1241
rect -29 -1309 29 -1275
rect -29 -1343 -17 -1309
rect 17 -1343 29 -1309
rect -29 -1377 29 -1343
rect -29 -1411 -17 -1377
rect 17 -1411 29 -1377
rect -29 -1445 29 -1411
rect -29 -1479 -17 -1445
rect 17 -1479 29 -1445
rect -29 -1513 29 -1479
rect -29 -1547 -17 -1513
rect 17 -1547 29 -1513
rect -29 -1581 29 -1547
rect -29 -1615 -17 -1581
rect 17 -1615 29 -1581
rect -29 -1649 29 -1615
rect -29 -1683 -17 -1649
rect 17 -1683 29 -1649
rect -29 -1717 29 -1683
rect -29 -1751 -17 -1717
rect 17 -1751 29 -1717
rect -29 -1785 29 -1751
rect -29 -1819 -17 -1785
rect 17 -1819 29 -1785
rect -29 -1853 29 -1819
rect -29 -1887 -17 -1853
rect 17 -1887 29 -1853
rect -29 -1900 29 -1887
rect 69 1887 127 1900
rect 69 1853 81 1887
rect 115 1853 127 1887
rect 69 1819 127 1853
rect 69 1785 81 1819
rect 115 1785 127 1819
rect 69 1751 127 1785
rect 69 1717 81 1751
rect 115 1717 127 1751
rect 69 1683 127 1717
rect 69 1649 81 1683
rect 115 1649 127 1683
rect 69 1615 127 1649
rect 69 1581 81 1615
rect 115 1581 127 1615
rect 69 1547 127 1581
rect 69 1513 81 1547
rect 115 1513 127 1547
rect 69 1479 127 1513
rect 69 1445 81 1479
rect 115 1445 127 1479
rect 69 1411 127 1445
rect 69 1377 81 1411
rect 115 1377 127 1411
rect 69 1343 127 1377
rect 69 1309 81 1343
rect 115 1309 127 1343
rect 69 1275 127 1309
rect 69 1241 81 1275
rect 115 1241 127 1275
rect 69 1207 127 1241
rect 69 1173 81 1207
rect 115 1173 127 1207
rect 69 1139 127 1173
rect 69 1105 81 1139
rect 115 1105 127 1139
rect 69 1071 127 1105
rect 69 1037 81 1071
rect 115 1037 127 1071
rect 69 1003 127 1037
rect 69 969 81 1003
rect 115 969 127 1003
rect 69 935 127 969
rect 69 901 81 935
rect 115 901 127 935
rect 69 867 127 901
rect 69 833 81 867
rect 115 833 127 867
rect 69 799 127 833
rect 69 765 81 799
rect 115 765 127 799
rect 69 731 127 765
rect 69 697 81 731
rect 115 697 127 731
rect 69 663 127 697
rect 69 629 81 663
rect 115 629 127 663
rect 69 595 127 629
rect 69 561 81 595
rect 115 561 127 595
rect 69 527 127 561
rect 69 493 81 527
rect 115 493 127 527
rect 69 459 127 493
rect 69 425 81 459
rect 115 425 127 459
rect 69 391 127 425
rect 69 357 81 391
rect 115 357 127 391
rect 69 323 127 357
rect 69 289 81 323
rect 115 289 127 323
rect 69 255 127 289
rect 69 221 81 255
rect 115 221 127 255
rect 69 187 127 221
rect 69 153 81 187
rect 115 153 127 187
rect 69 119 127 153
rect 69 85 81 119
rect 115 85 127 119
rect 69 51 127 85
rect 69 17 81 51
rect 115 17 127 51
rect 69 -17 127 17
rect 69 -51 81 -17
rect 115 -51 127 -17
rect 69 -85 127 -51
rect 69 -119 81 -85
rect 115 -119 127 -85
rect 69 -153 127 -119
rect 69 -187 81 -153
rect 115 -187 127 -153
rect 69 -221 127 -187
rect 69 -255 81 -221
rect 115 -255 127 -221
rect 69 -289 127 -255
rect 69 -323 81 -289
rect 115 -323 127 -289
rect 69 -357 127 -323
rect 69 -391 81 -357
rect 115 -391 127 -357
rect 69 -425 127 -391
rect 69 -459 81 -425
rect 115 -459 127 -425
rect 69 -493 127 -459
rect 69 -527 81 -493
rect 115 -527 127 -493
rect 69 -561 127 -527
rect 69 -595 81 -561
rect 115 -595 127 -561
rect 69 -629 127 -595
rect 69 -663 81 -629
rect 115 -663 127 -629
rect 69 -697 127 -663
rect 69 -731 81 -697
rect 115 -731 127 -697
rect 69 -765 127 -731
rect 69 -799 81 -765
rect 115 -799 127 -765
rect 69 -833 127 -799
rect 69 -867 81 -833
rect 115 -867 127 -833
rect 69 -901 127 -867
rect 69 -935 81 -901
rect 115 -935 127 -901
rect 69 -969 127 -935
rect 69 -1003 81 -969
rect 115 -1003 127 -969
rect 69 -1037 127 -1003
rect 69 -1071 81 -1037
rect 115 -1071 127 -1037
rect 69 -1105 127 -1071
rect 69 -1139 81 -1105
rect 115 -1139 127 -1105
rect 69 -1173 127 -1139
rect 69 -1207 81 -1173
rect 115 -1207 127 -1173
rect 69 -1241 127 -1207
rect 69 -1275 81 -1241
rect 115 -1275 127 -1241
rect 69 -1309 127 -1275
rect 69 -1343 81 -1309
rect 115 -1343 127 -1309
rect 69 -1377 127 -1343
rect 69 -1411 81 -1377
rect 115 -1411 127 -1377
rect 69 -1445 127 -1411
rect 69 -1479 81 -1445
rect 115 -1479 127 -1445
rect 69 -1513 127 -1479
rect 69 -1547 81 -1513
rect 115 -1547 127 -1513
rect 69 -1581 127 -1547
rect 69 -1615 81 -1581
rect 115 -1615 127 -1581
rect 69 -1649 127 -1615
rect 69 -1683 81 -1649
rect 115 -1683 127 -1649
rect 69 -1717 127 -1683
rect 69 -1751 81 -1717
rect 115 -1751 127 -1717
rect 69 -1785 127 -1751
rect 69 -1819 81 -1785
rect 115 -1819 127 -1785
rect 69 -1853 127 -1819
rect 69 -1887 81 -1853
rect 115 -1887 127 -1853
rect 69 -1900 127 -1887
rect 167 1887 225 1900
rect 167 1853 179 1887
rect 213 1853 225 1887
rect 167 1819 225 1853
rect 167 1785 179 1819
rect 213 1785 225 1819
rect 167 1751 225 1785
rect 167 1717 179 1751
rect 213 1717 225 1751
rect 167 1683 225 1717
rect 167 1649 179 1683
rect 213 1649 225 1683
rect 167 1615 225 1649
rect 167 1581 179 1615
rect 213 1581 225 1615
rect 167 1547 225 1581
rect 167 1513 179 1547
rect 213 1513 225 1547
rect 167 1479 225 1513
rect 167 1445 179 1479
rect 213 1445 225 1479
rect 167 1411 225 1445
rect 167 1377 179 1411
rect 213 1377 225 1411
rect 167 1343 225 1377
rect 167 1309 179 1343
rect 213 1309 225 1343
rect 167 1275 225 1309
rect 167 1241 179 1275
rect 213 1241 225 1275
rect 167 1207 225 1241
rect 167 1173 179 1207
rect 213 1173 225 1207
rect 167 1139 225 1173
rect 167 1105 179 1139
rect 213 1105 225 1139
rect 167 1071 225 1105
rect 167 1037 179 1071
rect 213 1037 225 1071
rect 167 1003 225 1037
rect 167 969 179 1003
rect 213 969 225 1003
rect 167 935 225 969
rect 167 901 179 935
rect 213 901 225 935
rect 167 867 225 901
rect 167 833 179 867
rect 213 833 225 867
rect 167 799 225 833
rect 167 765 179 799
rect 213 765 225 799
rect 167 731 225 765
rect 167 697 179 731
rect 213 697 225 731
rect 167 663 225 697
rect 167 629 179 663
rect 213 629 225 663
rect 167 595 225 629
rect 167 561 179 595
rect 213 561 225 595
rect 167 527 225 561
rect 167 493 179 527
rect 213 493 225 527
rect 167 459 225 493
rect 167 425 179 459
rect 213 425 225 459
rect 167 391 225 425
rect 167 357 179 391
rect 213 357 225 391
rect 167 323 225 357
rect 167 289 179 323
rect 213 289 225 323
rect 167 255 225 289
rect 167 221 179 255
rect 213 221 225 255
rect 167 187 225 221
rect 167 153 179 187
rect 213 153 225 187
rect 167 119 225 153
rect 167 85 179 119
rect 213 85 225 119
rect 167 51 225 85
rect 167 17 179 51
rect 213 17 225 51
rect 167 -17 225 17
rect 167 -51 179 -17
rect 213 -51 225 -17
rect 167 -85 225 -51
rect 167 -119 179 -85
rect 213 -119 225 -85
rect 167 -153 225 -119
rect 167 -187 179 -153
rect 213 -187 225 -153
rect 167 -221 225 -187
rect 167 -255 179 -221
rect 213 -255 225 -221
rect 167 -289 225 -255
rect 167 -323 179 -289
rect 213 -323 225 -289
rect 167 -357 225 -323
rect 167 -391 179 -357
rect 213 -391 225 -357
rect 167 -425 225 -391
rect 167 -459 179 -425
rect 213 -459 225 -425
rect 167 -493 225 -459
rect 167 -527 179 -493
rect 213 -527 225 -493
rect 167 -561 225 -527
rect 167 -595 179 -561
rect 213 -595 225 -561
rect 167 -629 225 -595
rect 167 -663 179 -629
rect 213 -663 225 -629
rect 167 -697 225 -663
rect 167 -731 179 -697
rect 213 -731 225 -697
rect 167 -765 225 -731
rect 167 -799 179 -765
rect 213 -799 225 -765
rect 167 -833 225 -799
rect 167 -867 179 -833
rect 213 -867 225 -833
rect 167 -901 225 -867
rect 167 -935 179 -901
rect 213 -935 225 -901
rect 167 -969 225 -935
rect 167 -1003 179 -969
rect 213 -1003 225 -969
rect 167 -1037 225 -1003
rect 167 -1071 179 -1037
rect 213 -1071 225 -1037
rect 167 -1105 225 -1071
rect 167 -1139 179 -1105
rect 213 -1139 225 -1105
rect 167 -1173 225 -1139
rect 167 -1207 179 -1173
rect 213 -1207 225 -1173
rect 167 -1241 225 -1207
rect 167 -1275 179 -1241
rect 213 -1275 225 -1241
rect 167 -1309 225 -1275
rect 167 -1343 179 -1309
rect 213 -1343 225 -1309
rect 167 -1377 225 -1343
rect 167 -1411 179 -1377
rect 213 -1411 225 -1377
rect 167 -1445 225 -1411
rect 167 -1479 179 -1445
rect 213 -1479 225 -1445
rect 167 -1513 225 -1479
rect 167 -1547 179 -1513
rect 213 -1547 225 -1513
rect 167 -1581 225 -1547
rect 167 -1615 179 -1581
rect 213 -1615 225 -1581
rect 167 -1649 225 -1615
rect 167 -1683 179 -1649
rect 213 -1683 225 -1649
rect 167 -1717 225 -1683
rect 167 -1751 179 -1717
rect 213 -1751 225 -1717
rect 167 -1785 225 -1751
rect 167 -1819 179 -1785
rect 213 -1819 225 -1785
rect 167 -1853 225 -1819
rect 167 -1887 179 -1853
rect 213 -1887 225 -1853
rect 167 -1900 225 -1887
<< pdiffc >>
rect -213 1853 -179 1887
rect -213 1785 -179 1819
rect -213 1717 -179 1751
rect -213 1649 -179 1683
rect -213 1581 -179 1615
rect -213 1513 -179 1547
rect -213 1445 -179 1479
rect -213 1377 -179 1411
rect -213 1309 -179 1343
rect -213 1241 -179 1275
rect -213 1173 -179 1207
rect -213 1105 -179 1139
rect -213 1037 -179 1071
rect -213 969 -179 1003
rect -213 901 -179 935
rect -213 833 -179 867
rect -213 765 -179 799
rect -213 697 -179 731
rect -213 629 -179 663
rect -213 561 -179 595
rect -213 493 -179 527
rect -213 425 -179 459
rect -213 357 -179 391
rect -213 289 -179 323
rect -213 221 -179 255
rect -213 153 -179 187
rect -213 85 -179 119
rect -213 17 -179 51
rect -213 -51 -179 -17
rect -213 -119 -179 -85
rect -213 -187 -179 -153
rect -213 -255 -179 -221
rect -213 -323 -179 -289
rect -213 -391 -179 -357
rect -213 -459 -179 -425
rect -213 -527 -179 -493
rect -213 -595 -179 -561
rect -213 -663 -179 -629
rect -213 -731 -179 -697
rect -213 -799 -179 -765
rect -213 -867 -179 -833
rect -213 -935 -179 -901
rect -213 -1003 -179 -969
rect -213 -1071 -179 -1037
rect -213 -1139 -179 -1105
rect -213 -1207 -179 -1173
rect -213 -1275 -179 -1241
rect -213 -1343 -179 -1309
rect -213 -1411 -179 -1377
rect -213 -1479 -179 -1445
rect -213 -1547 -179 -1513
rect -213 -1615 -179 -1581
rect -213 -1683 -179 -1649
rect -213 -1751 -179 -1717
rect -213 -1819 -179 -1785
rect -213 -1887 -179 -1853
rect -115 1853 -81 1887
rect -115 1785 -81 1819
rect -115 1717 -81 1751
rect -115 1649 -81 1683
rect -115 1581 -81 1615
rect -115 1513 -81 1547
rect -115 1445 -81 1479
rect -115 1377 -81 1411
rect -115 1309 -81 1343
rect -115 1241 -81 1275
rect -115 1173 -81 1207
rect -115 1105 -81 1139
rect -115 1037 -81 1071
rect -115 969 -81 1003
rect -115 901 -81 935
rect -115 833 -81 867
rect -115 765 -81 799
rect -115 697 -81 731
rect -115 629 -81 663
rect -115 561 -81 595
rect -115 493 -81 527
rect -115 425 -81 459
rect -115 357 -81 391
rect -115 289 -81 323
rect -115 221 -81 255
rect -115 153 -81 187
rect -115 85 -81 119
rect -115 17 -81 51
rect -115 -51 -81 -17
rect -115 -119 -81 -85
rect -115 -187 -81 -153
rect -115 -255 -81 -221
rect -115 -323 -81 -289
rect -115 -391 -81 -357
rect -115 -459 -81 -425
rect -115 -527 -81 -493
rect -115 -595 -81 -561
rect -115 -663 -81 -629
rect -115 -731 -81 -697
rect -115 -799 -81 -765
rect -115 -867 -81 -833
rect -115 -935 -81 -901
rect -115 -1003 -81 -969
rect -115 -1071 -81 -1037
rect -115 -1139 -81 -1105
rect -115 -1207 -81 -1173
rect -115 -1275 -81 -1241
rect -115 -1343 -81 -1309
rect -115 -1411 -81 -1377
rect -115 -1479 -81 -1445
rect -115 -1547 -81 -1513
rect -115 -1615 -81 -1581
rect -115 -1683 -81 -1649
rect -115 -1751 -81 -1717
rect -115 -1819 -81 -1785
rect -115 -1887 -81 -1853
rect -17 1853 17 1887
rect -17 1785 17 1819
rect -17 1717 17 1751
rect -17 1649 17 1683
rect -17 1581 17 1615
rect -17 1513 17 1547
rect -17 1445 17 1479
rect -17 1377 17 1411
rect -17 1309 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1139
rect -17 1037 17 1071
rect -17 969 17 1003
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1003 17 -969
rect -17 -1071 17 -1037
rect -17 -1139 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1309
rect -17 -1411 17 -1377
rect -17 -1479 17 -1445
rect -17 -1547 17 -1513
rect -17 -1615 17 -1581
rect -17 -1683 17 -1649
rect -17 -1751 17 -1717
rect -17 -1819 17 -1785
rect -17 -1887 17 -1853
rect 81 1853 115 1887
rect 81 1785 115 1819
rect 81 1717 115 1751
rect 81 1649 115 1683
rect 81 1581 115 1615
rect 81 1513 115 1547
rect 81 1445 115 1479
rect 81 1377 115 1411
rect 81 1309 115 1343
rect 81 1241 115 1275
rect 81 1173 115 1207
rect 81 1105 115 1139
rect 81 1037 115 1071
rect 81 969 115 1003
rect 81 901 115 935
rect 81 833 115 867
rect 81 765 115 799
rect 81 697 115 731
rect 81 629 115 663
rect 81 561 115 595
rect 81 493 115 527
rect 81 425 115 459
rect 81 357 115 391
rect 81 289 115 323
rect 81 221 115 255
rect 81 153 115 187
rect 81 85 115 119
rect 81 17 115 51
rect 81 -51 115 -17
rect 81 -119 115 -85
rect 81 -187 115 -153
rect 81 -255 115 -221
rect 81 -323 115 -289
rect 81 -391 115 -357
rect 81 -459 115 -425
rect 81 -527 115 -493
rect 81 -595 115 -561
rect 81 -663 115 -629
rect 81 -731 115 -697
rect 81 -799 115 -765
rect 81 -867 115 -833
rect 81 -935 115 -901
rect 81 -1003 115 -969
rect 81 -1071 115 -1037
rect 81 -1139 115 -1105
rect 81 -1207 115 -1173
rect 81 -1275 115 -1241
rect 81 -1343 115 -1309
rect 81 -1411 115 -1377
rect 81 -1479 115 -1445
rect 81 -1547 115 -1513
rect 81 -1615 115 -1581
rect 81 -1683 115 -1649
rect 81 -1751 115 -1717
rect 81 -1819 115 -1785
rect 81 -1887 115 -1853
rect 179 1853 213 1887
rect 179 1785 213 1819
rect 179 1717 213 1751
rect 179 1649 213 1683
rect 179 1581 213 1615
rect 179 1513 213 1547
rect 179 1445 213 1479
rect 179 1377 213 1411
rect 179 1309 213 1343
rect 179 1241 213 1275
rect 179 1173 213 1207
rect 179 1105 213 1139
rect 179 1037 213 1071
rect 179 969 213 1003
rect 179 901 213 935
rect 179 833 213 867
rect 179 765 213 799
rect 179 697 213 731
rect 179 629 213 663
rect 179 561 213 595
rect 179 493 213 527
rect 179 425 213 459
rect 179 357 213 391
rect 179 289 213 323
rect 179 221 213 255
rect 179 153 213 187
rect 179 85 213 119
rect 179 17 213 51
rect 179 -51 213 -17
rect 179 -119 213 -85
rect 179 -187 213 -153
rect 179 -255 213 -221
rect 179 -323 213 -289
rect 179 -391 213 -357
rect 179 -459 213 -425
rect 179 -527 213 -493
rect 179 -595 213 -561
rect 179 -663 213 -629
rect 179 -731 213 -697
rect 179 -799 213 -765
rect 179 -867 213 -833
rect 179 -935 213 -901
rect 179 -1003 213 -969
rect 179 -1071 213 -1037
rect 179 -1139 213 -1105
rect 179 -1207 213 -1173
rect 179 -1275 213 -1241
rect 179 -1343 213 -1309
rect 179 -1411 213 -1377
rect 179 -1479 213 -1445
rect 179 -1547 213 -1513
rect 179 -1615 213 -1581
rect 179 -1683 213 -1649
rect 179 -1751 213 -1717
rect 179 -1819 213 -1785
rect 179 -1887 213 -1853
<< nsubdiff >>
rect -327 2049 -221 2083
rect -187 2049 -153 2083
rect -119 2049 -85 2083
rect -51 2049 -17 2083
rect 17 2049 51 2083
rect 85 2049 119 2083
rect 153 2049 187 2083
rect 221 2049 327 2083
rect -327 1955 -293 2049
rect 293 1955 327 2049
rect -327 1887 -293 1921
rect -327 1819 -293 1853
rect -327 1751 -293 1785
rect -327 1683 -293 1717
rect -327 1615 -293 1649
rect -327 1547 -293 1581
rect -327 1479 -293 1513
rect -327 1411 -293 1445
rect -327 1343 -293 1377
rect -327 1275 -293 1309
rect -327 1207 -293 1241
rect -327 1139 -293 1173
rect -327 1071 -293 1105
rect -327 1003 -293 1037
rect -327 935 -293 969
rect -327 867 -293 901
rect -327 799 -293 833
rect -327 731 -293 765
rect -327 663 -293 697
rect -327 595 -293 629
rect -327 527 -293 561
rect -327 459 -293 493
rect -327 391 -293 425
rect -327 323 -293 357
rect -327 255 -293 289
rect -327 187 -293 221
rect -327 119 -293 153
rect -327 51 -293 85
rect -327 -17 -293 17
rect -327 -85 -293 -51
rect -327 -153 -293 -119
rect -327 -221 -293 -187
rect -327 -289 -293 -255
rect -327 -357 -293 -323
rect -327 -425 -293 -391
rect -327 -493 -293 -459
rect -327 -561 -293 -527
rect -327 -629 -293 -595
rect -327 -697 -293 -663
rect -327 -765 -293 -731
rect -327 -833 -293 -799
rect -327 -901 -293 -867
rect -327 -969 -293 -935
rect -327 -1037 -293 -1003
rect -327 -1105 -293 -1071
rect -327 -1173 -293 -1139
rect -327 -1241 -293 -1207
rect -327 -1309 -293 -1275
rect -327 -1377 -293 -1343
rect -327 -1445 -293 -1411
rect -327 -1513 -293 -1479
rect -327 -1581 -293 -1547
rect -327 -1649 -293 -1615
rect -327 -1717 -293 -1683
rect -327 -1785 -293 -1751
rect -327 -1853 -293 -1819
rect -327 -1921 -293 -1887
rect 293 1887 327 1921
rect 293 1819 327 1853
rect 293 1751 327 1785
rect 293 1683 327 1717
rect 293 1615 327 1649
rect 293 1547 327 1581
rect 293 1479 327 1513
rect 293 1411 327 1445
rect 293 1343 327 1377
rect 293 1275 327 1309
rect 293 1207 327 1241
rect 293 1139 327 1173
rect 293 1071 327 1105
rect 293 1003 327 1037
rect 293 935 327 969
rect 293 867 327 901
rect 293 799 327 833
rect 293 731 327 765
rect 293 663 327 697
rect 293 595 327 629
rect 293 527 327 561
rect 293 459 327 493
rect 293 391 327 425
rect 293 323 327 357
rect 293 255 327 289
rect 293 187 327 221
rect 293 119 327 153
rect 293 51 327 85
rect 293 -17 327 17
rect 293 -85 327 -51
rect 293 -153 327 -119
rect 293 -221 327 -187
rect 293 -289 327 -255
rect 293 -357 327 -323
rect 293 -425 327 -391
rect 293 -493 327 -459
rect 293 -561 327 -527
rect 293 -629 327 -595
rect 293 -697 327 -663
rect 293 -765 327 -731
rect 293 -833 327 -799
rect 293 -901 327 -867
rect 293 -969 327 -935
rect 293 -1037 327 -1003
rect 293 -1105 327 -1071
rect 293 -1173 327 -1139
rect 293 -1241 327 -1207
rect 293 -1309 327 -1275
rect 293 -1377 327 -1343
rect 293 -1445 327 -1411
rect 293 -1513 327 -1479
rect 293 -1581 327 -1547
rect 293 -1649 327 -1615
rect 293 -1717 327 -1683
rect 293 -1785 327 -1751
rect 293 -1853 327 -1819
rect 293 -1921 327 -1887
rect -327 -2049 -293 -1955
rect 293 -2049 327 -1955
rect -327 -2083 -221 -2049
rect -187 -2083 -153 -2049
rect -119 -2083 -85 -2049
rect -51 -2083 -17 -2049
rect 17 -2083 51 -2049
rect 85 -2083 119 -2049
rect 153 -2083 187 -2049
rect 221 -2083 327 -2049
<< nsubdiffcont >>
rect -221 2049 -187 2083
rect -153 2049 -119 2083
rect -85 2049 -51 2083
rect -17 2049 17 2083
rect 51 2049 85 2083
rect 119 2049 153 2083
rect 187 2049 221 2083
rect -327 1921 -293 1955
rect 293 1921 327 1955
rect -327 1853 -293 1887
rect -327 1785 -293 1819
rect -327 1717 -293 1751
rect -327 1649 -293 1683
rect -327 1581 -293 1615
rect -327 1513 -293 1547
rect -327 1445 -293 1479
rect -327 1377 -293 1411
rect -327 1309 -293 1343
rect -327 1241 -293 1275
rect -327 1173 -293 1207
rect -327 1105 -293 1139
rect -327 1037 -293 1071
rect -327 969 -293 1003
rect -327 901 -293 935
rect -327 833 -293 867
rect -327 765 -293 799
rect -327 697 -293 731
rect -327 629 -293 663
rect -327 561 -293 595
rect -327 493 -293 527
rect -327 425 -293 459
rect -327 357 -293 391
rect -327 289 -293 323
rect -327 221 -293 255
rect -327 153 -293 187
rect -327 85 -293 119
rect -327 17 -293 51
rect -327 -51 -293 -17
rect -327 -119 -293 -85
rect -327 -187 -293 -153
rect -327 -255 -293 -221
rect -327 -323 -293 -289
rect -327 -391 -293 -357
rect -327 -459 -293 -425
rect -327 -527 -293 -493
rect -327 -595 -293 -561
rect -327 -663 -293 -629
rect -327 -731 -293 -697
rect -327 -799 -293 -765
rect -327 -867 -293 -833
rect -327 -935 -293 -901
rect -327 -1003 -293 -969
rect -327 -1071 -293 -1037
rect -327 -1139 -293 -1105
rect -327 -1207 -293 -1173
rect -327 -1275 -293 -1241
rect -327 -1343 -293 -1309
rect -327 -1411 -293 -1377
rect -327 -1479 -293 -1445
rect -327 -1547 -293 -1513
rect -327 -1615 -293 -1581
rect -327 -1683 -293 -1649
rect -327 -1751 -293 -1717
rect -327 -1819 -293 -1785
rect -327 -1887 -293 -1853
rect 293 1853 327 1887
rect 293 1785 327 1819
rect 293 1717 327 1751
rect 293 1649 327 1683
rect 293 1581 327 1615
rect 293 1513 327 1547
rect 293 1445 327 1479
rect 293 1377 327 1411
rect 293 1309 327 1343
rect 293 1241 327 1275
rect 293 1173 327 1207
rect 293 1105 327 1139
rect 293 1037 327 1071
rect 293 969 327 1003
rect 293 901 327 935
rect 293 833 327 867
rect 293 765 327 799
rect 293 697 327 731
rect 293 629 327 663
rect 293 561 327 595
rect 293 493 327 527
rect 293 425 327 459
rect 293 357 327 391
rect 293 289 327 323
rect 293 221 327 255
rect 293 153 327 187
rect 293 85 327 119
rect 293 17 327 51
rect 293 -51 327 -17
rect 293 -119 327 -85
rect 293 -187 327 -153
rect 293 -255 327 -221
rect 293 -323 327 -289
rect 293 -391 327 -357
rect 293 -459 327 -425
rect 293 -527 327 -493
rect 293 -595 327 -561
rect 293 -663 327 -629
rect 293 -731 327 -697
rect 293 -799 327 -765
rect 293 -867 327 -833
rect 293 -935 327 -901
rect 293 -1003 327 -969
rect 293 -1071 327 -1037
rect 293 -1139 327 -1105
rect 293 -1207 327 -1173
rect 293 -1275 327 -1241
rect 293 -1343 327 -1309
rect 293 -1411 327 -1377
rect 293 -1479 327 -1445
rect 293 -1547 327 -1513
rect 293 -1615 327 -1581
rect 293 -1683 327 -1649
rect 293 -1751 327 -1717
rect 293 -1819 327 -1785
rect 293 -1887 327 -1853
rect -327 -1955 -293 -1921
rect 293 -1955 327 -1921
rect -221 -2083 -187 -2049
rect -153 -2083 -119 -2049
rect -85 -2083 -51 -2049
rect -17 -2083 17 -2049
rect 51 -2083 85 -2049
rect 119 -2083 153 -2049
rect 187 -2083 221 -2049
<< poly >>
rect -82 1981 -16 1997
rect -82 1947 -66 1981
rect -32 1947 -16 1981
rect -82 1931 -16 1947
rect 114 1981 180 1997
rect 114 1947 130 1981
rect 164 1947 180 1981
rect 114 1931 180 1947
rect -167 1900 -127 1926
rect -69 1900 -29 1931
rect 29 1900 69 1926
rect 127 1900 167 1931
rect -167 -1931 -127 -1900
rect -69 -1926 -29 -1900
rect 29 -1931 69 -1900
rect 127 -1926 167 -1900
rect -180 -1947 -114 -1931
rect -180 -1981 -164 -1947
rect -130 -1981 -114 -1947
rect -180 -1997 -114 -1981
rect 16 -1947 82 -1931
rect 16 -1981 32 -1947
rect 66 -1981 82 -1947
rect 16 -1997 82 -1981
<< polycont >>
rect -66 1947 -32 1981
rect 130 1947 164 1981
rect -164 -1981 -130 -1947
rect 32 -1981 66 -1947
<< locali >>
rect -327 2049 -221 2083
rect -187 2049 -153 2083
rect -119 2049 -85 2083
rect -51 2049 -17 2083
rect 17 2049 51 2083
rect 85 2049 119 2083
rect 153 2049 187 2083
rect 221 2049 327 2083
rect -327 1955 -293 2049
rect -82 1947 -66 1981
rect -32 1947 -16 1981
rect 114 1947 130 1981
rect 164 1947 180 1981
rect 293 1955 327 2049
rect -327 1887 -293 1921
rect -327 1819 -293 1853
rect -327 1751 -293 1785
rect -327 1683 -293 1717
rect -327 1615 -293 1649
rect -327 1547 -293 1581
rect -327 1479 -293 1513
rect -327 1411 -293 1445
rect -327 1343 -293 1377
rect -327 1275 -293 1309
rect -327 1207 -293 1241
rect -327 1139 -293 1173
rect -327 1071 -293 1105
rect -327 1003 -293 1037
rect -327 935 -293 969
rect -327 867 -293 901
rect -327 799 -293 833
rect -327 731 -293 765
rect -327 663 -293 697
rect -327 595 -293 629
rect -327 527 -293 561
rect -327 459 -293 493
rect -327 391 -293 425
rect -327 323 -293 357
rect -327 255 -293 289
rect -327 187 -293 221
rect -327 119 -293 153
rect -327 51 -293 85
rect -327 -17 -293 17
rect -327 -85 -293 -51
rect -327 -153 -293 -119
rect -327 -221 -293 -187
rect -327 -289 -293 -255
rect -327 -357 -293 -323
rect -327 -425 -293 -391
rect -327 -493 -293 -459
rect -327 -561 -293 -527
rect -327 -629 -293 -595
rect -327 -697 -293 -663
rect -327 -765 -293 -731
rect -327 -833 -293 -799
rect -327 -901 -293 -867
rect -327 -969 -293 -935
rect -327 -1037 -293 -1003
rect -327 -1105 -293 -1071
rect -327 -1173 -293 -1139
rect -327 -1241 -293 -1207
rect -327 -1309 -293 -1275
rect -327 -1377 -293 -1343
rect -327 -1445 -293 -1411
rect -327 -1513 -293 -1479
rect -327 -1581 -293 -1547
rect -327 -1649 -293 -1615
rect -327 -1717 -293 -1683
rect -327 -1785 -293 -1751
rect -327 -1853 -293 -1819
rect -327 -1921 -293 -1887
rect -213 1887 -179 1904
rect -213 1781 -179 1785
rect -213 1709 -179 1717
rect -213 1637 -179 1649
rect -213 1565 -179 1581
rect -213 1493 -179 1513
rect -213 1421 -179 1445
rect -213 1349 -179 1377
rect -213 1277 -179 1309
rect -213 1207 -179 1241
rect -213 1139 -179 1171
rect -213 1071 -179 1099
rect -213 1003 -179 1027
rect -213 935 -179 955
rect -213 867 -179 883
rect -213 799 -179 811
rect -213 731 -179 739
rect -213 663 -179 667
rect -213 557 -179 561
rect -213 485 -179 493
rect -213 413 -179 425
rect -213 341 -179 357
rect -213 269 -179 289
rect -213 197 -179 221
rect -213 125 -179 153
rect -213 53 -179 85
rect -213 -17 -179 17
rect -213 -85 -179 -53
rect -213 -153 -179 -125
rect -213 -221 -179 -197
rect -213 -289 -179 -269
rect -213 -357 -179 -341
rect -213 -425 -179 -413
rect -213 -493 -179 -485
rect -213 -561 -179 -557
rect -213 -667 -179 -663
rect -213 -739 -179 -731
rect -213 -811 -179 -799
rect -213 -883 -179 -867
rect -213 -955 -179 -935
rect -213 -1027 -179 -1003
rect -213 -1099 -179 -1071
rect -213 -1171 -179 -1139
rect -213 -1241 -179 -1207
rect -213 -1309 -179 -1277
rect -213 -1377 -179 -1349
rect -213 -1445 -179 -1421
rect -213 -1513 -179 -1493
rect -213 -1581 -179 -1565
rect -213 -1649 -179 -1637
rect -213 -1717 -179 -1709
rect -213 -1785 -179 -1781
rect -213 -1904 -179 -1887
rect -115 1887 -81 1904
rect -115 1781 -81 1785
rect -115 1709 -81 1717
rect -115 1637 -81 1649
rect -115 1565 -81 1581
rect -115 1493 -81 1513
rect -115 1421 -81 1445
rect -115 1349 -81 1377
rect -115 1277 -81 1309
rect -115 1207 -81 1241
rect -115 1139 -81 1171
rect -115 1071 -81 1099
rect -115 1003 -81 1027
rect -115 935 -81 955
rect -115 867 -81 883
rect -115 799 -81 811
rect -115 731 -81 739
rect -115 663 -81 667
rect -115 557 -81 561
rect -115 485 -81 493
rect -115 413 -81 425
rect -115 341 -81 357
rect -115 269 -81 289
rect -115 197 -81 221
rect -115 125 -81 153
rect -115 53 -81 85
rect -115 -17 -81 17
rect -115 -85 -81 -53
rect -115 -153 -81 -125
rect -115 -221 -81 -197
rect -115 -289 -81 -269
rect -115 -357 -81 -341
rect -115 -425 -81 -413
rect -115 -493 -81 -485
rect -115 -561 -81 -557
rect -115 -667 -81 -663
rect -115 -739 -81 -731
rect -115 -811 -81 -799
rect -115 -883 -81 -867
rect -115 -955 -81 -935
rect -115 -1027 -81 -1003
rect -115 -1099 -81 -1071
rect -115 -1171 -81 -1139
rect -115 -1241 -81 -1207
rect -115 -1309 -81 -1277
rect -115 -1377 -81 -1349
rect -115 -1445 -81 -1421
rect -115 -1513 -81 -1493
rect -115 -1581 -81 -1565
rect -115 -1649 -81 -1637
rect -115 -1717 -81 -1709
rect -115 -1785 -81 -1781
rect -115 -1904 -81 -1887
rect -17 1887 17 1904
rect -17 1781 17 1785
rect -17 1709 17 1717
rect -17 1637 17 1649
rect -17 1565 17 1581
rect -17 1493 17 1513
rect -17 1421 17 1445
rect -17 1349 17 1377
rect -17 1277 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1171
rect -17 1071 17 1099
rect -17 1003 17 1027
rect -17 935 17 955
rect -17 867 17 883
rect -17 799 17 811
rect -17 731 17 739
rect -17 663 17 667
rect -17 557 17 561
rect -17 485 17 493
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -493 17 -485
rect -17 -561 17 -557
rect -17 -667 17 -663
rect -17 -739 17 -731
rect -17 -811 17 -799
rect -17 -883 17 -867
rect -17 -955 17 -935
rect -17 -1027 17 -1003
rect -17 -1099 17 -1071
rect -17 -1171 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1277
rect -17 -1377 17 -1349
rect -17 -1445 17 -1421
rect -17 -1513 17 -1493
rect -17 -1581 17 -1565
rect -17 -1649 17 -1637
rect -17 -1717 17 -1709
rect -17 -1785 17 -1781
rect -17 -1904 17 -1887
rect 81 1887 115 1904
rect 81 1781 115 1785
rect 81 1709 115 1717
rect 81 1637 115 1649
rect 81 1565 115 1581
rect 81 1493 115 1513
rect 81 1421 115 1445
rect 81 1349 115 1377
rect 81 1277 115 1309
rect 81 1207 115 1241
rect 81 1139 115 1171
rect 81 1071 115 1099
rect 81 1003 115 1027
rect 81 935 115 955
rect 81 867 115 883
rect 81 799 115 811
rect 81 731 115 739
rect 81 663 115 667
rect 81 557 115 561
rect 81 485 115 493
rect 81 413 115 425
rect 81 341 115 357
rect 81 269 115 289
rect 81 197 115 221
rect 81 125 115 153
rect 81 53 115 85
rect 81 -17 115 17
rect 81 -85 115 -53
rect 81 -153 115 -125
rect 81 -221 115 -197
rect 81 -289 115 -269
rect 81 -357 115 -341
rect 81 -425 115 -413
rect 81 -493 115 -485
rect 81 -561 115 -557
rect 81 -667 115 -663
rect 81 -739 115 -731
rect 81 -811 115 -799
rect 81 -883 115 -867
rect 81 -955 115 -935
rect 81 -1027 115 -1003
rect 81 -1099 115 -1071
rect 81 -1171 115 -1139
rect 81 -1241 115 -1207
rect 81 -1309 115 -1277
rect 81 -1377 115 -1349
rect 81 -1445 115 -1421
rect 81 -1513 115 -1493
rect 81 -1581 115 -1565
rect 81 -1649 115 -1637
rect 81 -1717 115 -1709
rect 81 -1785 115 -1781
rect 81 -1904 115 -1887
rect 179 1887 213 1904
rect 179 1781 213 1785
rect 179 1709 213 1717
rect 179 1637 213 1649
rect 179 1565 213 1581
rect 179 1493 213 1513
rect 179 1421 213 1445
rect 179 1349 213 1377
rect 179 1277 213 1309
rect 179 1207 213 1241
rect 179 1139 213 1171
rect 179 1071 213 1099
rect 179 1003 213 1027
rect 179 935 213 955
rect 179 867 213 883
rect 179 799 213 811
rect 179 731 213 739
rect 179 663 213 667
rect 179 557 213 561
rect 179 485 213 493
rect 179 413 213 425
rect 179 341 213 357
rect 179 269 213 289
rect 179 197 213 221
rect 179 125 213 153
rect 179 53 213 85
rect 179 -17 213 17
rect 179 -85 213 -53
rect 179 -153 213 -125
rect 179 -221 213 -197
rect 179 -289 213 -269
rect 179 -357 213 -341
rect 179 -425 213 -413
rect 179 -493 213 -485
rect 179 -561 213 -557
rect 179 -667 213 -663
rect 179 -739 213 -731
rect 179 -811 213 -799
rect 179 -883 213 -867
rect 179 -955 213 -935
rect 179 -1027 213 -1003
rect 179 -1099 213 -1071
rect 179 -1171 213 -1139
rect 179 -1241 213 -1207
rect 179 -1309 213 -1277
rect 179 -1377 213 -1349
rect 179 -1445 213 -1421
rect 179 -1513 213 -1493
rect 179 -1581 213 -1565
rect 179 -1649 213 -1637
rect 179 -1717 213 -1709
rect 179 -1785 213 -1781
rect 179 -1904 213 -1887
rect 293 1887 327 1921
rect 293 1819 327 1853
rect 293 1751 327 1785
rect 293 1683 327 1717
rect 293 1615 327 1649
rect 293 1547 327 1581
rect 293 1479 327 1513
rect 293 1411 327 1445
rect 293 1343 327 1377
rect 293 1275 327 1309
rect 293 1207 327 1241
rect 293 1139 327 1173
rect 293 1071 327 1105
rect 293 1003 327 1037
rect 293 935 327 969
rect 293 867 327 901
rect 293 799 327 833
rect 293 731 327 765
rect 293 663 327 697
rect 293 595 327 629
rect 293 527 327 561
rect 293 459 327 493
rect 293 391 327 425
rect 293 323 327 357
rect 293 255 327 289
rect 293 187 327 221
rect 293 119 327 153
rect 293 51 327 85
rect 293 -17 327 17
rect 293 -85 327 -51
rect 293 -153 327 -119
rect 293 -221 327 -187
rect 293 -289 327 -255
rect 293 -357 327 -323
rect 293 -425 327 -391
rect 293 -493 327 -459
rect 293 -561 327 -527
rect 293 -629 327 -595
rect 293 -697 327 -663
rect 293 -765 327 -731
rect 293 -833 327 -799
rect 293 -901 327 -867
rect 293 -969 327 -935
rect 293 -1037 327 -1003
rect 293 -1105 327 -1071
rect 293 -1173 327 -1139
rect 293 -1241 327 -1207
rect 293 -1309 327 -1275
rect 293 -1377 327 -1343
rect 293 -1445 327 -1411
rect 293 -1513 327 -1479
rect 293 -1581 327 -1547
rect 293 -1649 327 -1615
rect 293 -1717 327 -1683
rect 293 -1785 327 -1751
rect 293 -1853 327 -1819
rect 293 -1921 327 -1887
rect -327 -2049 -293 -1955
rect -180 -1981 -164 -1947
rect -130 -1981 -114 -1947
rect 16 -1981 32 -1947
rect 66 -1981 82 -1947
rect 293 -2049 327 -1955
rect -327 -2083 -221 -2049
rect -187 -2083 -153 -2049
rect -119 -2083 -85 -2049
rect -51 -2083 -17 -2049
rect 17 -2083 51 -2049
rect 85 -2083 119 -2049
rect 153 -2083 187 -2049
rect 221 -2083 327 -2049
<< viali >>
rect -66 1947 -32 1981
rect 130 1947 164 1981
rect -213 1819 -179 1853
rect -213 1751 -179 1781
rect -213 1747 -179 1751
rect -213 1683 -179 1709
rect -213 1675 -179 1683
rect -213 1615 -179 1637
rect -213 1603 -179 1615
rect -213 1547 -179 1565
rect -213 1531 -179 1547
rect -213 1479 -179 1493
rect -213 1459 -179 1479
rect -213 1411 -179 1421
rect -213 1387 -179 1411
rect -213 1343 -179 1349
rect -213 1315 -179 1343
rect -213 1275 -179 1277
rect -213 1243 -179 1275
rect -213 1173 -179 1205
rect -213 1171 -179 1173
rect -213 1105 -179 1133
rect -213 1099 -179 1105
rect -213 1037 -179 1061
rect -213 1027 -179 1037
rect -213 969 -179 989
rect -213 955 -179 969
rect -213 901 -179 917
rect -213 883 -179 901
rect -213 833 -179 845
rect -213 811 -179 833
rect -213 765 -179 773
rect -213 739 -179 765
rect -213 697 -179 701
rect -213 667 -179 697
rect -213 595 -179 629
rect -213 527 -179 557
rect -213 523 -179 527
rect -213 459 -179 485
rect -213 451 -179 459
rect -213 391 -179 413
rect -213 379 -179 391
rect -213 323 -179 341
rect -213 307 -179 323
rect -213 255 -179 269
rect -213 235 -179 255
rect -213 187 -179 197
rect -213 163 -179 187
rect -213 119 -179 125
rect -213 91 -179 119
rect -213 51 -179 53
rect -213 19 -179 51
rect -213 -51 -179 -19
rect -213 -53 -179 -51
rect -213 -119 -179 -91
rect -213 -125 -179 -119
rect -213 -187 -179 -163
rect -213 -197 -179 -187
rect -213 -255 -179 -235
rect -213 -269 -179 -255
rect -213 -323 -179 -307
rect -213 -341 -179 -323
rect -213 -391 -179 -379
rect -213 -413 -179 -391
rect -213 -459 -179 -451
rect -213 -485 -179 -459
rect -213 -527 -179 -523
rect -213 -557 -179 -527
rect -213 -629 -179 -595
rect -213 -697 -179 -667
rect -213 -701 -179 -697
rect -213 -765 -179 -739
rect -213 -773 -179 -765
rect -213 -833 -179 -811
rect -213 -845 -179 -833
rect -213 -901 -179 -883
rect -213 -917 -179 -901
rect -213 -969 -179 -955
rect -213 -989 -179 -969
rect -213 -1037 -179 -1027
rect -213 -1061 -179 -1037
rect -213 -1105 -179 -1099
rect -213 -1133 -179 -1105
rect -213 -1173 -179 -1171
rect -213 -1205 -179 -1173
rect -213 -1275 -179 -1243
rect -213 -1277 -179 -1275
rect -213 -1343 -179 -1315
rect -213 -1349 -179 -1343
rect -213 -1411 -179 -1387
rect -213 -1421 -179 -1411
rect -213 -1479 -179 -1459
rect -213 -1493 -179 -1479
rect -213 -1547 -179 -1531
rect -213 -1565 -179 -1547
rect -213 -1615 -179 -1603
rect -213 -1637 -179 -1615
rect -213 -1683 -179 -1675
rect -213 -1709 -179 -1683
rect -213 -1751 -179 -1747
rect -213 -1781 -179 -1751
rect -213 -1853 -179 -1819
rect -115 1819 -81 1853
rect -115 1751 -81 1781
rect -115 1747 -81 1751
rect -115 1683 -81 1709
rect -115 1675 -81 1683
rect -115 1615 -81 1637
rect -115 1603 -81 1615
rect -115 1547 -81 1565
rect -115 1531 -81 1547
rect -115 1479 -81 1493
rect -115 1459 -81 1479
rect -115 1411 -81 1421
rect -115 1387 -81 1411
rect -115 1343 -81 1349
rect -115 1315 -81 1343
rect -115 1275 -81 1277
rect -115 1243 -81 1275
rect -115 1173 -81 1205
rect -115 1171 -81 1173
rect -115 1105 -81 1133
rect -115 1099 -81 1105
rect -115 1037 -81 1061
rect -115 1027 -81 1037
rect -115 969 -81 989
rect -115 955 -81 969
rect -115 901 -81 917
rect -115 883 -81 901
rect -115 833 -81 845
rect -115 811 -81 833
rect -115 765 -81 773
rect -115 739 -81 765
rect -115 697 -81 701
rect -115 667 -81 697
rect -115 595 -81 629
rect -115 527 -81 557
rect -115 523 -81 527
rect -115 459 -81 485
rect -115 451 -81 459
rect -115 391 -81 413
rect -115 379 -81 391
rect -115 323 -81 341
rect -115 307 -81 323
rect -115 255 -81 269
rect -115 235 -81 255
rect -115 187 -81 197
rect -115 163 -81 187
rect -115 119 -81 125
rect -115 91 -81 119
rect -115 51 -81 53
rect -115 19 -81 51
rect -115 -51 -81 -19
rect -115 -53 -81 -51
rect -115 -119 -81 -91
rect -115 -125 -81 -119
rect -115 -187 -81 -163
rect -115 -197 -81 -187
rect -115 -255 -81 -235
rect -115 -269 -81 -255
rect -115 -323 -81 -307
rect -115 -341 -81 -323
rect -115 -391 -81 -379
rect -115 -413 -81 -391
rect -115 -459 -81 -451
rect -115 -485 -81 -459
rect -115 -527 -81 -523
rect -115 -557 -81 -527
rect -115 -629 -81 -595
rect -115 -697 -81 -667
rect -115 -701 -81 -697
rect -115 -765 -81 -739
rect -115 -773 -81 -765
rect -115 -833 -81 -811
rect -115 -845 -81 -833
rect -115 -901 -81 -883
rect -115 -917 -81 -901
rect -115 -969 -81 -955
rect -115 -989 -81 -969
rect -115 -1037 -81 -1027
rect -115 -1061 -81 -1037
rect -115 -1105 -81 -1099
rect -115 -1133 -81 -1105
rect -115 -1173 -81 -1171
rect -115 -1205 -81 -1173
rect -115 -1275 -81 -1243
rect -115 -1277 -81 -1275
rect -115 -1343 -81 -1315
rect -115 -1349 -81 -1343
rect -115 -1411 -81 -1387
rect -115 -1421 -81 -1411
rect -115 -1479 -81 -1459
rect -115 -1493 -81 -1479
rect -115 -1547 -81 -1531
rect -115 -1565 -81 -1547
rect -115 -1615 -81 -1603
rect -115 -1637 -81 -1615
rect -115 -1683 -81 -1675
rect -115 -1709 -81 -1683
rect -115 -1751 -81 -1747
rect -115 -1781 -81 -1751
rect -115 -1853 -81 -1819
rect -17 1819 17 1853
rect -17 1751 17 1781
rect -17 1747 17 1751
rect -17 1683 17 1709
rect -17 1675 17 1683
rect -17 1615 17 1637
rect -17 1603 17 1615
rect -17 1547 17 1565
rect -17 1531 17 1547
rect -17 1479 17 1493
rect -17 1459 17 1479
rect -17 1411 17 1421
rect -17 1387 17 1411
rect -17 1343 17 1349
rect -17 1315 17 1343
rect -17 1275 17 1277
rect -17 1243 17 1275
rect -17 1173 17 1205
rect -17 1171 17 1173
rect -17 1105 17 1133
rect -17 1099 17 1105
rect -17 1037 17 1061
rect -17 1027 17 1037
rect -17 969 17 989
rect -17 955 17 969
rect -17 901 17 917
rect -17 883 17 901
rect -17 833 17 845
rect -17 811 17 833
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect -17 -833 17 -811
rect -17 -845 17 -833
rect -17 -901 17 -883
rect -17 -917 17 -901
rect -17 -969 17 -955
rect -17 -989 17 -969
rect -17 -1037 17 -1027
rect -17 -1061 17 -1037
rect -17 -1105 17 -1099
rect -17 -1133 17 -1105
rect -17 -1173 17 -1171
rect -17 -1205 17 -1173
rect -17 -1275 17 -1243
rect -17 -1277 17 -1275
rect -17 -1343 17 -1315
rect -17 -1349 17 -1343
rect -17 -1411 17 -1387
rect -17 -1421 17 -1411
rect -17 -1479 17 -1459
rect -17 -1493 17 -1479
rect -17 -1547 17 -1531
rect -17 -1565 17 -1547
rect -17 -1615 17 -1603
rect -17 -1637 17 -1615
rect -17 -1683 17 -1675
rect -17 -1709 17 -1683
rect -17 -1751 17 -1747
rect -17 -1781 17 -1751
rect -17 -1853 17 -1819
rect 81 1819 115 1853
rect 81 1751 115 1781
rect 81 1747 115 1751
rect 81 1683 115 1709
rect 81 1675 115 1683
rect 81 1615 115 1637
rect 81 1603 115 1615
rect 81 1547 115 1565
rect 81 1531 115 1547
rect 81 1479 115 1493
rect 81 1459 115 1479
rect 81 1411 115 1421
rect 81 1387 115 1411
rect 81 1343 115 1349
rect 81 1315 115 1343
rect 81 1275 115 1277
rect 81 1243 115 1275
rect 81 1173 115 1205
rect 81 1171 115 1173
rect 81 1105 115 1133
rect 81 1099 115 1105
rect 81 1037 115 1061
rect 81 1027 115 1037
rect 81 969 115 989
rect 81 955 115 969
rect 81 901 115 917
rect 81 883 115 901
rect 81 833 115 845
rect 81 811 115 833
rect 81 765 115 773
rect 81 739 115 765
rect 81 697 115 701
rect 81 667 115 697
rect 81 595 115 629
rect 81 527 115 557
rect 81 523 115 527
rect 81 459 115 485
rect 81 451 115 459
rect 81 391 115 413
rect 81 379 115 391
rect 81 323 115 341
rect 81 307 115 323
rect 81 255 115 269
rect 81 235 115 255
rect 81 187 115 197
rect 81 163 115 187
rect 81 119 115 125
rect 81 91 115 119
rect 81 51 115 53
rect 81 19 115 51
rect 81 -51 115 -19
rect 81 -53 115 -51
rect 81 -119 115 -91
rect 81 -125 115 -119
rect 81 -187 115 -163
rect 81 -197 115 -187
rect 81 -255 115 -235
rect 81 -269 115 -255
rect 81 -323 115 -307
rect 81 -341 115 -323
rect 81 -391 115 -379
rect 81 -413 115 -391
rect 81 -459 115 -451
rect 81 -485 115 -459
rect 81 -527 115 -523
rect 81 -557 115 -527
rect 81 -629 115 -595
rect 81 -697 115 -667
rect 81 -701 115 -697
rect 81 -765 115 -739
rect 81 -773 115 -765
rect 81 -833 115 -811
rect 81 -845 115 -833
rect 81 -901 115 -883
rect 81 -917 115 -901
rect 81 -969 115 -955
rect 81 -989 115 -969
rect 81 -1037 115 -1027
rect 81 -1061 115 -1037
rect 81 -1105 115 -1099
rect 81 -1133 115 -1105
rect 81 -1173 115 -1171
rect 81 -1205 115 -1173
rect 81 -1275 115 -1243
rect 81 -1277 115 -1275
rect 81 -1343 115 -1315
rect 81 -1349 115 -1343
rect 81 -1411 115 -1387
rect 81 -1421 115 -1411
rect 81 -1479 115 -1459
rect 81 -1493 115 -1479
rect 81 -1547 115 -1531
rect 81 -1565 115 -1547
rect 81 -1615 115 -1603
rect 81 -1637 115 -1615
rect 81 -1683 115 -1675
rect 81 -1709 115 -1683
rect 81 -1751 115 -1747
rect 81 -1781 115 -1751
rect 81 -1853 115 -1819
rect 179 1819 213 1853
rect 179 1751 213 1781
rect 179 1747 213 1751
rect 179 1683 213 1709
rect 179 1675 213 1683
rect 179 1615 213 1637
rect 179 1603 213 1615
rect 179 1547 213 1565
rect 179 1531 213 1547
rect 179 1479 213 1493
rect 179 1459 213 1479
rect 179 1411 213 1421
rect 179 1387 213 1411
rect 179 1343 213 1349
rect 179 1315 213 1343
rect 179 1275 213 1277
rect 179 1243 213 1275
rect 179 1173 213 1205
rect 179 1171 213 1173
rect 179 1105 213 1133
rect 179 1099 213 1105
rect 179 1037 213 1061
rect 179 1027 213 1037
rect 179 969 213 989
rect 179 955 213 969
rect 179 901 213 917
rect 179 883 213 901
rect 179 833 213 845
rect 179 811 213 833
rect 179 765 213 773
rect 179 739 213 765
rect 179 697 213 701
rect 179 667 213 697
rect 179 595 213 629
rect 179 527 213 557
rect 179 523 213 527
rect 179 459 213 485
rect 179 451 213 459
rect 179 391 213 413
rect 179 379 213 391
rect 179 323 213 341
rect 179 307 213 323
rect 179 255 213 269
rect 179 235 213 255
rect 179 187 213 197
rect 179 163 213 187
rect 179 119 213 125
rect 179 91 213 119
rect 179 51 213 53
rect 179 19 213 51
rect 179 -51 213 -19
rect 179 -53 213 -51
rect 179 -119 213 -91
rect 179 -125 213 -119
rect 179 -187 213 -163
rect 179 -197 213 -187
rect 179 -255 213 -235
rect 179 -269 213 -255
rect 179 -323 213 -307
rect 179 -341 213 -323
rect 179 -391 213 -379
rect 179 -413 213 -391
rect 179 -459 213 -451
rect 179 -485 213 -459
rect 179 -527 213 -523
rect 179 -557 213 -527
rect 179 -629 213 -595
rect 179 -697 213 -667
rect 179 -701 213 -697
rect 179 -765 213 -739
rect 179 -773 213 -765
rect 179 -833 213 -811
rect 179 -845 213 -833
rect 179 -901 213 -883
rect 179 -917 213 -901
rect 179 -969 213 -955
rect 179 -989 213 -969
rect 179 -1037 213 -1027
rect 179 -1061 213 -1037
rect 179 -1105 213 -1099
rect 179 -1133 213 -1105
rect 179 -1173 213 -1171
rect 179 -1205 213 -1173
rect 179 -1275 213 -1243
rect 179 -1277 213 -1275
rect 179 -1343 213 -1315
rect 179 -1349 213 -1343
rect 179 -1411 213 -1387
rect 179 -1421 213 -1411
rect 179 -1479 213 -1459
rect 179 -1493 213 -1479
rect 179 -1547 213 -1531
rect 179 -1565 213 -1547
rect 179 -1615 213 -1603
rect 179 -1637 213 -1615
rect 179 -1683 213 -1675
rect 179 -1709 213 -1683
rect 179 -1751 213 -1747
rect 179 -1781 213 -1751
rect 179 -1853 213 -1819
rect -164 -1981 -130 -1947
rect 32 -1981 66 -1947
<< metal1 >>
rect -78 1981 -20 1987
rect -78 1947 -66 1981
rect -32 1947 -20 1981
rect -78 1941 -20 1947
rect 118 1981 176 1987
rect 118 1947 130 1981
rect 164 1947 176 1981
rect 118 1941 176 1947
rect -219 1853 -173 1900
rect -219 1819 -213 1853
rect -179 1819 -173 1853
rect -219 1781 -173 1819
rect -219 1747 -213 1781
rect -179 1747 -173 1781
rect -219 1709 -173 1747
rect -219 1675 -213 1709
rect -179 1675 -173 1709
rect -219 1637 -173 1675
rect -219 1603 -213 1637
rect -179 1603 -173 1637
rect -219 1565 -173 1603
rect -219 1531 -213 1565
rect -179 1531 -173 1565
rect -219 1493 -173 1531
rect -219 1459 -213 1493
rect -179 1459 -173 1493
rect -219 1421 -173 1459
rect -219 1387 -213 1421
rect -179 1387 -173 1421
rect -219 1349 -173 1387
rect -219 1315 -213 1349
rect -179 1315 -173 1349
rect -219 1277 -173 1315
rect -219 1243 -213 1277
rect -179 1243 -173 1277
rect -219 1205 -173 1243
rect -219 1171 -213 1205
rect -179 1171 -173 1205
rect -219 1133 -173 1171
rect -219 1099 -213 1133
rect -179 1099 -173 1133
rect -219 1061 -173 1099
rect -219 1027 -213 1061
rect -179 1027 -173 1061
rect -219 989 -173 1027
rect -219 955 -213 989
rect -179 955 -173 989
rect -219 917 -173 955
rect -219 883 -213 917
rect -179 883 -173 917
rect -219 845 -173 883
rect -219 811 -213 845
rect -179 811 -173 845
rect -219 773 -173 811
rect -219 739 -213 773
rect -179 739 -173 773
rect -219 701 -173 739
rect -219 667 -213 701
rect -179 667 -173 701
rect -219 629 -173 667
rect -219 595 -213 629
rect -179 595 -173 629
rect -219 557 -173 595
rect -219 523 -213 557
rect -179 523 -173 557
rect -219 485 -173 523
rect -219 451 -213 485
rect -179 451 -173 485
rect -219 413 -173 451
rect -219 379 -213 413
rect -179 379 -173 413
rect -219 341 -173 379
rect -219 307 -213 341
rect -179 307 -173 341
rect -219 269 -173 307
rect -219 235 -213 269
rect -179 235 -173 269
rect -219 197 -173 235
rect -219 163 -213 197
rect -179 163 -173 197
rect -219 125 -173 163
rect -219 91 -213 125
rect -179 91 -173 125
rect -219 53 -173 91
rect -219 19 -213 53
rect -179 19 -173 53
rect -219 -19 -173 19
rect -219 -53 -213 -19
rect -179 -53 -173 -19
rect -219 -91 -173 -53
rect -219 -125 -213 -91
rect -179 -125 -173 -91
rect -219 -163 -173 -125
rect -219 -197 -213 -163
rect -179 -197 -173 -163
rect -219 -235 -173 -197
rect -219 -269 -213 -235
rect -179 -269 -173 -235
rect -219 -307 -173 -269
rect -219 -341 -213 -307
rect -179 -341 -173 -307
rect -219 -379 -173 -341
rect -219 -413 -213 -379
rect -179 -413 -173 -379
rect -219 -451 -173 -413
rect -219 -485 -213 -451
rect -179 -485 -173 -451
rect -219 -523 -173 -485
rect -219 -557 -213 -523
rect -179 -557 -173 -523
rect -219 -595 -173 -557
rect -219 -629 -213 -595
rect -179 -629 -173 -595
rect -219 -667 -173 -629
rect -219 -701 -213 -667
rect -179 -701 -173 -667
rect -219 -739 -173 -701
rect -219 -773 -213 -739
rect -179 -773 -173 -739
rect -219 -811 -173 -773
rect -219 -845 -213 -811
rect -179 -845 -173 -811
rect -219 -883 -173 -845
rect -219 -917 -213 -883
rect -179 -917 -173 -883
rect -219 -955 -173 -917
rect -219 -989 -213 -955
rect -179 -989 -173 -955
rect -219 -1027 -173 -989
rect -219 -1061 -213 -1027
rect -179 -1061 -173 -1027
rect -219 -1099 -173 -1061
rect -219 -1133 -213 -1099
rect -179 -1133 -173 -1099
rect -219 -1171 -173 -1133
rect -219 -1205 -213 -1171
rect -179 -1205 -173 -1171
rect -219 -1243 -173 -1205
rect -219 -1277 -213 -1243
rect -179 -1277 -173 -1243
rect -219 -1315 -173 -1277
rect -219 -1349 -213 -1315
rect -179 -1349 -173 -1315
rect -219 -1387 -173 -1349
rect -219 -1421 -213 -1387
rect -179 -1421 -173 -1387
rect -219 -1459 -173 -1421
rect -219 -1493 -213 -1459
rect -179 -1493 -173 -1459
rect -219 -1531 -173 -1493
rect -219 -1565 -213 -1531
rect -179 -1565 -173 -1531
rect -219 -1603 -173 -1565
rect -219 -1637 -213 -1603
rect -179 -1637 -173 -1603
rect -219 -1675 -173 -1637
rect -219 -1709 -213 -1675
rect -179 -1709 -173 -1675
rect -219 -1747 -173 -1709
rect -219 -1781 -213 -1747
rect -179 -1781 -173 -1747
rect -219 -1819 -173 -1781
rect -219 -1853 -213 -1819
rect -179 -1853 -173 -1819
rect -219 -1900 -173 -1853
rect -121 1853 -75 1900
rect -121 1819 -115 1853
rect -81 1819 -75 1853
rect -121 1781 -75 1819
rect -121 1747 -115 1781
rect -81 1747 -75 1781
rect -121 1709 -75 1747
rect -121 1675 -115 1709
rect -81 1675 -75 1709
rect -121 1637 -75 1675
rect -121 1603 -115 1637
rect -81 1603 -75 1637
rect -121 1565 -75 1603
rect -121 1531 -115 1565
rect -81 1531 -75 1565
rect -121 1493 -75 1531
rect -121 1459 -115 1493
rect -81 1459 -75 1493
rect -121 1421 -75 1459
rect -121 1387 -115 1421
rect -81 1387 -75 1421
rect -121 1349 -75 1387
rect -121 1315 -115 1349
rect -81 1315 -75 1349
rect -121 1277 -75 1315
rect -121 1243 -115 1277
rect -81 1243 -75 1277
rect -121 1205 -75 1243
rect -121 1171 -115 1205
rect -81 1171 -75 1205
rect -121 1133 -75 1171
rect -121 1099 -115 1133
rect -81 1099 -75 1133
rect -121 1061 -75 1099
rect -121 1027 -115 1061
rect -81 1027 -75 1061
rect -121 989 -75 1027
rect -121 955 -115 989
rect -81 955 -75 989
rect -121 917 -75 955
rect -121 883 -115 917
rect -81 883 -75 917
rect -121 845 -75 883
rect -121 811 -115 845
rect -81 811 -75 845
rect -121 773 -75 811
rect -121 739 -115 773
rect -81 739 -75 773
rect -121 701 -75 739
rect -121 667 -115 701
rect -81 667 -75 701
rect -121 629 -75 667
rect -121 595 -115 629
rect -81 595 -75 629
rect -121 557 -75 595
rect -121 523 -115 557
rect -81 523 -75 557
rect -121 485 -75 523
rect -121 451 -115 485
rect -81 451 -75 485
rect -121 413 -75 451
rect -121 379 -115 413
rect -81 379 -75 413
rect -121 341 -75 379
rect -121 307 -115 341
rect -81 307 -75 341
rect -121 269 -75 307
rect -121 235 -115 269
rect -81 235 -75 269
rect -121 197 -75 235
rect -121 163 -115 197
rect -81 163 -75 197
rect -121 125 -75 163
rect -121 91 -115 125
rect -81 91 -75 125
rect -121 53 -75 91
rect -121 19 -115 53
rect -81 19 -75 53
rect -121 -19 -75 19
rect -121 -53 -115 -19
rect -81 -53 -75 -19
rect -121 -91 -75 -53
rect -121 -125 -115 -91
rect -81 -125 -75 -91
rect -121 -163 -75 -125
rect -121 -197 -115 -163
rect -81 -197 -75 -163
rect -121 -235 -75 -197
rect -121 -269 -115 -235
rect -81 -269 -75 -235
rect -121 -307 -75 -269
rect -121 -341 -115 -307
rect -81 -341 -75 -307
rect -121 -379 -75 -341
rect -121 -413 -115 -379
rect -81 -413 -75 -379
rect -121 -451 -75 -413
rect -121 -485 -115 -451
rect -81 -485 -75 -451
rect -121 -523 -75 -485
rect -121 -557 -115 -523
rect -81 -557 -75 -523
rect -121 -595 -75 -557
rect -121 -629 -115 -595
rect -81 -629 -75 -595
rect -121 -667 -75 -629
rect -121 -701 -115 -667
rect -81 -701 -75 -667
rect -121 -739 -75 -701
rect -121 -773 -115 -739
rect -81 -773 -75 -739
rect -121 -811 -75 -773
rect -121 -845 -115 -811
rect -81 -845 -75 -811
rect -121 -883 -75 -845
rect -121 -917 -115 -883
rect -81 -917 -75 -883
rect -121 -955 -75 -917
rect -121 -989 -115 -955
rect -81 -989 -75 -955
rect -121 -1027 -75 -989
rect -121 -1061 -115 -1027
rect -81 -1061 -75 -1027
rect -121 -1099 -75 -1061
rect -121 -1133 -115 -1099
rect -81 -1133 -75 -1099
rect -121 -1171 -75 -1133
rect -121 -1205 -115 -1171
rect -81 -1205 -75 -1171
rect -121 -1243 -75 -1205
rect -121 -1277 -115 -1243
rect -81 -1277 -75 -1243
rect -121 -1315 -75 -1277
rect -121 -1349 -115 -1315
rect -81 -1349 -75 -1315
rect -121 -1387 -75 -1349
rect -121 -1421 -115 -1387
rect -81 -1421 -75 -1387
rect -121 -1459 -75 -1421
rect -121 -1493 -115 -1459
rect -81 -1493 -75 -1459
rect -121 -1531 -75 -1493
rect -121 -1565 -115 -1531
rect -81 -1565 -75 -1531
rect -121 -1603 -75 -1565
rect -121 -1637 -115 -1603
rect -81 -1637 -75 -1603
rect -121 -1675 -75 -1637
rect -121 -1709 -115 -1675
rect -81 -1709 -75 -1675
rect -121 -1747 -75 -1709
rect -121 -1781 -115 -1747
rect -81 -1781 -75 -1747
rect -121 -1819 -75 -1781
rect -121 -1853 -115 -1819
rect -81 -1853 -75 -1819
rect -121 -1900 -75 -1853
rect -23 1853 23 1900
rect -23 1819 -17 1853
rect 17 1819 23 1853
rect -23 1781 23 1819
rect -23 1747 -17 1781
rect 17 1747 23 1781
rect -23 1709 23 1747
rect -23 1675 -17 1709
rect 17 1675 23 1709
rect -23 1637 23 1675
rect -23 1603 -17 1637
rect 17 1603 23 1637
rect -23 1565 23 1603
rect -23 1531 -17 1565
rect 17 1531 23 1565
rect -23 1493 23 1531
rect -23 1459 -17 1493
rect 17 1459 23 1493
rect -23 1421 23 1459
rect -23 1387 -17 1421
rect 17 1387 23 1421
rect -23 1349 23 1387
rect -23 1315 -17 1349
rect 17 1315 23 1349
rect -23 1277 23 1315
rect -23 1243 -17 1277
rect 17 1243 23 1277
rect -23 1205 23 1243
rect -23 1171 -17 1205
rect 17 1171 23 1205
rect -23 1133 23 1171
rect -23 1099 -17 1133
rect 17 1099 23 1133
rect -23 1061 23 1099
rect -23 1027 -17 1061
rect 17 1027 23 1061
rect -23 989 23 1027
rect -23 955 -17 989
rect 17 955 23 989
rect -23 917 23 955
rect -23 883 -17 917
rect 17 883 23 917
rect -23 845 23 883
rect -23 811 -17 845
rect 17 811 23 845
rect -23 773 23 811
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -811 23 -773
rect -23 -845 -17 -811
rect 17 -845 23 -811
rect -23 -883 23 -845
rect -23 -917 -17 -883
rect 17 -917 23 -883
rect -23 -955 23 -917
rect -23 -989 -17 -955
rect 17 -989 23 -955
rect -23 -1027 23 -989
rect -23 -1061 -17 -1027
rect 17 -1061 23 -1027
rect -23 -1099 23 -1061
rect -23 -1133 -17 -1099
rect 17 -1133 23 -1099
rect -23 -1171 23 -1133
rect -23 -1205 -17 -1171
rect 17 -1205 23 -1171
rect -23 -1243 23 -1205
rect -23 -1277 -17 -1243
rect 17 -1277 23 -1243
rect -23 -1315 23 -1277
rect -23 -1349 -17 -1315
rect 17 -1349 23 -1315
rect -23 -1387 23 -1349
rect -23 -1421 -17 -1387
rect 17 -1421 23 -1387
rect -23 -1459 23 -1421
rect -23 -1493 -17 -1459
rect 17 -1493 23 -1459
rect -23 -1531 23 -1493
rect -23 -1565 -17 -1531
rect 17 -1565 23 -1531
rect -23 -1603 23 -1565
rect -23 -1637 -17 -1603
rect 17 -1637 23 -1603
rect -23 -1675 23 -1637
rect -23 -1709 -17 -1675
rect 17 -1709 23 -1675
rect -23 -1747 23 -1709
rect -23 -1781 -17 -1747
rect 17 -1781 23 -1747
rect -23 -1819 23 -1781
rect -23 -1853 -17 -1819
rect 17 -1853 23 -1819
rect -23 -1900 23 -1853
rect 75 1853 121 1900
rect 75 1819 81 1853
rect 115 1819 121 1853
rect 75 1781 121 1819
rect 75 1747 81 1781
rect 115 1747 121 1781
rect 75 1709 121 1747
rect 75 1675 81 1709
rect 115 1675 121 1709
rect 75 1637 121 1675
rect 75 1603 81 1637
rect 115 1603 121 1637
rect 75 1565 121 1603
rect 75 1531 81 1565
rect 115 1531 121 1565
rect 75 1493 121 1531
rect 75 1459 81 1493
rect 115 1459 121 1493
rect 75 1421 121 1459
rect 75 1387 81 1421
rect 115 1387 121 1421
rect 75 1349 121 1387
rect 75 1315 81 1349
rect 115 1315 121 1349
rect 75 1277 121 1315
rect 75 1243 81 1277
rect 115 1243 121 1277
rect 75 1205 121 1243
rect 75 1171 81 1205
rect 115 1171 121 1205
rect 75 1133 121 1171
rect 75 1099 81 1133
rect 115 1099 121 1133
rect 75 1061 121 1099
rect 75 1027 81 1061
rect 115 1027 121 1061
rect 75 989 121 1027
rect 75 955 81 989
rect 115 955 121 989
rect 75 917 121 955
rect 75 883 81 917
rect 115 883 121 917
rect 75 845 121 883
rect 75 811 81 845
rect 115 811 121 845
rect 75 773 121 811
rect 75 739 81 773
rect 115 739 121 773
rect 75 701 121 739
rect 75 667 81 701
rect 115 667 121 701
rect 75 629 121 667
rect 75 595 81 629
rect 115 595 121 629
rect 75 557 121 595
rect 75 523 81 557
rect 115 523 121 557
rect 75 485 121 523
rect 75 451 81 485
rect 115 451 121 485
rect 75 413 121 451
rect 75 379 81 413
rect 115 379 121 413
rect 75 341 121 379
rect 75 307 81 341
rect 115 307 121 341
rect 75 269 121 307
rect 75 235 81 269
rect 115 235 121 269
rect 75 197 121 235
rect 75 163 81 197
rect 115 163 121 197
rect 75 125 121 163
rect 75 91 81 125
rect 115 91 121 125
rect 75 53 121 91
rect 75 19 81 53
rect 115 19 121 53
rect 75 -19 121 19
rect 75 -53 81 -19
rect 115 -53 121 -19
rect 75 -91 121 -53
rect 75 -125 81 -91
rect 115 -125 121 -91
rect 75 -163 121 -125
rect 75 -197 81 -163
rect 115 -197 121 -163
rect 75 -235 121 -197
rect 75 -269 81 -235
rect 115 -269 121 -235
rect 75 -307 121 -269
rect 75 -341 81 -307
rect 115 -341 121 -307
rect 75 -379 121 -341
rect 75 -413 81 -379
rect 115 -413 121 -379
rect 75 -451 121 -413
rect 75 -485 81 -451
rect 115 -485 121 -451
rect 75 -523 121 -485
rect 75 -557 81 -523
rect 115 -557 121 -523
rect 75 -595 121 -557
rect 75 -629 81 -595
rect 115 -629 121 -595
rect 75 -667 121 -629
rect 75 -701 81 -667
rect 115 -701 121 -667
rect 75 -739 121 -701
rect 75 -773 81 -739
rect 115 -773 121 -739
rect 75 -811 121 -773
rect 75 -845 81 -811
rect 115 -845 121 -811
rect 75 -883 121 -845
rect 75 -917 81 -883
rect 115 -917 121 -883
rect 75 -955 121 -917
rect 75 -989 81 -955
rect 115 -989 121 -955
rect 75 -1027 121 -989
rect 75 -1061 81 -1027
rect 115 -1061 121 -1027
rect 75 -1099 121 -1061
rect 75 -1133 81 -1099
rect 115 -1133 121 -1099
rect 75 -1171 121 -1133
rect 75 -1205 81 -1171
rect 115 -1205 121 -1171
rect 75 -1243 121 -1205
rect 75 -1277 81 -1243
rect 115 -1277 121 -1243
rect 75 -1315 121 -1277
rect 75 -1349 81 -1315
rect 115 -1349 121 -1315
rect 75 -1387 121 -1349
rect 75 -1421 81 -1387
rect 115 -1421 121 -1387
rect 75 -1459 121 -1421
rect 75 -1493 81 -1459
rect 115 -1493 121 -1459
rect 75 -1531 121 -1493
rect 75 -1565 81 -1531
rect 115 -1565 121 -1531
rect 75 -1603 121 -1565
rect 75 -1637 81 -1603
rect 115 -1637 121 -1603
rect 75 -1675 121 -1637
rect 75 -1709 81 -1675
rect 115 -1709 121 -1675
rect 75 -1747 121 -1709
rect 75 -1781 81 -1747
rect 115 -1781 121 -1747
rect 75 -1819 121 -1781
rect 75 -1853 81 -1819
rect 115 -1853 121 -1819
rect 75 -1900 121 -1853
rect 173 1853 219 1900
rect 173 1819 179 1853
rect 213 1819 219 1853
rect 173 1781 219 1819
rect 173 1747 179 1781
rect 213 1747 219 1781
rect 173 1709 219 1747
rect 173 1675 179 1709
rect 213 1675 219 1709
rect 173 1637 219 1675
rect 173 1603 179 1637
rect 213 1603 219 1637
rect 173 1565 219 1603
rect 173 1531 179 1565
rect 213 1531 219 1565
rect 173 1493 219 1531
rect 173 1459 179 1493
rect 213 1459 219 1493
rect 173 1421 219 1459
rect 173 1387 179 1421
rect 213 1387 219 1421
rect 173 1349 219 1387
rect 173 1315 179 1349
rect 213 1315 219 1349
rect 173 1277 219 1315
rect 173 1243 179 1277
rect 213 1243 219 1277
rect 173 1205 219 1243
rect 173 1171 179 1205
rect 213 1171 219 1205
rect 173 1133 219 1171
rect 173 1099 179 1133
rect 213 1099 219 1133
rect 173 1061 219 1099
rect 173 1027 179 1061
rect 213 1027 219 1061
rect 173 989 219 1027
rect 173 955 179 989
rect 213 955 219 989
rect 173 917 219 955
rect 173 883 179 917
rect 213 883 219 917
rect 173 845 219 883
rect 173 811 179 845
rect 213 811 219 845
rect 173 773 219 811
rect 173 739 179 773
rect 213 739 219 773
rect 173 701 219 739
rect 173 667 179 701
rect 213 667 219 701
rect 173 629 219 667
rect 173 595 179 629
rect 213 595 219 629
rect 173 557 219 595
rect 173 523 179 557
rect 213 523 219 557
rect 173 485 219 523
rect 173 451 179 485
rect 213 451 219 485
rect 173 413 219 451
rect 173 379 179 413
rect 213 379 219 413
rect 173 341 219 379
rect 173 307 179 341
rect 213 307 219 341
rect 173 269 219 307
rect 173 235 179 269
rect 213 235 219 269
rect 173 197 219 235
rect 173 163 179 197
rect 213 163 219 197
rect 173 125 219 163
rect 173 91 179 125
rect 213 91 219 125
rect 173 53 219 91
rect 173 19 179 53
rect 213 19 219 53
rect 173 -19 219 19
rect 173 -53 179 -19
rect 213 -53 219 -19
rect 173 -91 219 -53
rect 173 -125 179 -91
rect 213 -125 219 -91
rect 173 -163 219 -125
rect 173 -197 179 -163
rect 213 -197 219 -163
rect 173 -235 219 -197
rect 173 -269 179 -235
rect 213 -269 219 -235
rect 173 -307 219 -269
rect 173 -341 179 -307
rect 213 -341 219 -307
rect 173 -379 219 -341
rect 173 -413 179 -379
rect 213 -413 219 -379
rect 173 -451 219 -413
rect 173 -485 179 -451
rect 213 -485 219 -451
rect 173 -523 219 -485
rect 173 -557 179 -523
rect 213 -557 219 -523
rect 173 -595 219 -557
rect 173 -629 179 -595
rect 213 -629 219 -595
rect 173 -667 219 -629
rect 173 -701 179 -667
rect 213 -701 219 -667
rect 173 -739 219 -701
rect 173 -773 179 -739
rect 213 -773 219 -739
rect 173 -811 219 -773
rect 173 -845 179 -811
rect 213 -845 219 -811
rect 173 -883 219 -845
rect 173 -917 179 -883
rect 213 -917 219 -883
rect 173 -955 219 -917
rect 173 -989 179 -955
rect 213 -989 219 -955
rect 173 -1027 219 -989
rect 173 -1061 179 -1027
rect 213 -1061 219 -1027
rect 173 -1099 219 -1061
rect 173 -1133 179 -1099
rect 213 -1133 219 -1099
rect 173 -1171 219 -1133
rect 173 -1205 179 -1171
rect 213 -1205 219 -1171
rect 173 -1243 219 -1205
rect 173 -1277 179 -1243
rect 213 -1277 219 -1243
rect 173 -1315 219 -1277
rect 173 -1349 179 -1315
rect 213 -1349 219 -1315
rect 173 -1387 219 -1349
rect 173 -1421 179 -1387
rect 213 -1421 219 -1387
rect 173 -1459 219 -1421
rect 173 -1493 179 -1459
rect 213 -1493 219 -1459
rect 173 -1531 219 -1493
rect 173 -1565 179 -1531
rect 213 -1565 219 -1531
rect 173 -1603 219 -1565
rect 173 -1637 179 -1603
rect 213 -1637 219 -1603
rect 173 -1675 219 -1637
rect 173 -1709 179 -1675
rect 213 -1709 219 -1675
rect 173 -1747 219 -1709
rect 173 -1781 179 -1747
rect 213 -1781 219 -1747
rect 173 -1819 219 -1781
rect 173 -1853 179 -1819
rect 213 -1853 219 -1819
rect 173 -1900 219 -1853
rect -176 -1947 -118 -1941
rect -176 -1981 -164 -1947
rect -130 -1981 -118 -1947
rect -176 -1987 -118 -1981
rect 20 -1947 78 -1941
rect 20 -1981 32 -1947
rect 66 -1981 78 -1947
rect 20 -1987 78 -1981
<< properties >>
string FIXED_BBOX -310 -2066 310 2066
<< end >>
