magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -246 -419 246 419
<< pmos >>
rect -50 -200 50 200
<< pdiff >>
rect -108 187 -50 200
rect -108 153 -96 187
rect -62 153 -50 187
rect -108 119 -50 153
rect -108 85 -96 119
rect -62 85 -50 119
rect -108 51 -50 85
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -85 -50 -51
rect -108 -119 -96 -85
rect -62 -119 -50 -85
rect -108 -153 -50 -119
rect -108 -187 -96 -153
rect -62 -187 -50 -153
rect -108 -200 -50 -187
rect 50 187 108 200
rect 50 153 62 187
rect 96 153 108 187
rect 50 119 108 153
rect 50 85 62 119
rect 96 85 108 119
rect 50 51 108 85
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -85 108 -51
rect 50 -119 62 -85
rect 96 -119 108 -85
rect 50 -153 108 -119
rect 50 -187 62 -153
rect 96 -187 108 -153
rect 50 -200 108 -187
<< pdiffc >>
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
<< nsubdiff >>
rect -210 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 210 383
rect -210 255 -176 349
rect -210 187 -176 221
rect 176 255 210 349
rect -210 119 -176 153
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect 176 187 210 221
rect 176 119 210 153
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect 176 -153 210 -119
rect -210 -349 -176 -255
rect 176 -221 210 -187
rect 176 -349 210 -255
rect -210 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 210 -349
<< nsubdiffcont >>
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect -210 221 -176 255
rect 176 221 210 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect -210 -255 -176 -221
rect 176 -255 210 -221
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
<< poly >>
rect -50 281 50 297
rect -50 247 -17 281
rect 17 247 50 281
rect -50 200 50 247
rect -50 -247 50 -200
rect -50 -281 -17 -247
rect 17 -281 50 -247
rect -50 -297 50 -281
<< polycont >>
rect -17 247 17 281
rect -17 -281 17 -247
<< locali >>
rect -210 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 210 383
rect -210 255 -176 349
rect -50 247 -17 281
rect 17 247 50 281
rect 176 255 210 349
rect -210 187 -176 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -96 187 -62 204
rect -96 119 -62 127
rect -96 51 -62 55
rect -96 -55 -62 -51
rect -96 -127 -62 -119
rect -96 -204 -62 -187
rect 62 187 96 204
rect 62 119 96 127
rect 62 51 96 55
rect 62 -55 96 -51
rect 62 -127 96 -119
rect 62 -204 96 -187
rect 176 187 210 221
rect 176 119 210 153
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect -210 -349 -176 -255
rect -50 -281 -17 -247
rect 17 -281 50 -247
rect 176 -349 210 -255
rect -210 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 210 -349
<< viali >>
rect -17 247 17 281
rect -96 153 -62 161
rect -96 127 -62 153
rect -96 85 -62 89
rect -96 55 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -55
rect -96 -89 -62 -85
rect -96 -153 -62 -127
rect -96 -161 -62 -153
rect 62 153 96 161
rect 62 127 96 153
rect 62 85 96 89
rect 62 55 96 85
rect 62 -17 96 17
rect 62 -85 96 -55
rect 62 -89 96 -85
rect 62 -153 96 -127
rect 62 -161 96 -153
rect -17 -281 17 -247
<< metal1 >>
rect -46 281 46 287
rect -46 247 -17 281
rect 17 247 46 281
rect -46 241 46 247
rect -102 161 -56 200
rect -102 127 -96 161
rect -62 127 -56 161
rect -102 89 -56 127
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -127 -56 -89
rect -102 -161 -96 -127
rect -62 -161 -56 -127
rect -102 -200 -56 -161
rect 56 161 102 200
rect 56 127 62 161
rect 96 127 102 161
rect 56 89 102 127
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -127 102 -89
rect 56 -161 62 -127
rect 96 -161 102 -127
rect 56 -200 102 -161
rect -46 -247 46 -241
rect -46 -281 -17 -247
rect 17 -281 46 -247
rect -46 -287 46 -281
<< properties >>
string FIXED_BBOX -193 -366 193 366
<< end >>
