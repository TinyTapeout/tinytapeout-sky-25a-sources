// Generated from: 20250915-070516_binTestAcc9760_seed230646_epochs100_2x4000_b256_lr30_interconnect.npz

module net (
    input  wire [253:0] in,
    output wire [3999:0] out,
    output wire [2549:0] categories
);
    wire [4000:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = in[137] & ~in[53]; 
    assign layer_0[1] = ~(in[98] ^ in[85]); 
    assign layer_0[2] = ~(in[117] | in[88]); 
    assign layer_0[3] = in[88] ^ in[197]; 
    assign layer_0[4] = ~in[168] | (in[168] & in[163]); 
    assign layer_0[5] = ~(in[39] ^ in[134]); 
    assign layer_0[6] = ~(in[38] ^ in[66]); 
    assign layer_0[7] = ~(in[147] ^ in[149]); 
    assign layer_0[8] = ~(in[186] | in[63]); 
    assign layer_0[9] = in[131]; 
    assign layer_0[10] = ~(in[219] ^ in[251]); 
    assign layer_0[11] = in[138] & ~in[164]; 
    assign layer_0[12] = ~(in[101] | in[197]); 
    assign layer_0[13] = ~(in[138] | in[124]); 
    assign layer_0[14] = ~(in[153] ^ in[114]); 
    assign layer_0[15] = in[59]; 
    assign layer_0[16] = ~(in[242] | in[250]); 
    assign layer_0[17] = in[102] & ~in[113]; 
    assign layer_0[18] = ~(in[132] ^ in[166]); 
    assign layer_0[19] = in[250] ^ in[164]; 
    assign layer_0[20] = ~(in[103] ^ in[54]); 
    assign layer_0[21] = in[9]; 
    assign layer_0[22] = ~(in[219] | in[58]); 
    assign layer_0[23] = in[217] | in[77]; 
    assign layer_0[24] = in[154] & ~in[173]; 
    assign layer_0[25] = in[115]; 
    assign layer_0[26] = in[116] & ~in[137]; 
    assign layer_0[27] = ~in[87] | (in[87] & in[52]); 
    assign layer_0[28] = in[71] & ~in[151]; 
    assign layer_0[29] = ~(in[55] ^ in[197]); 
    assign layer_0[30] = in[103] ^ in[107]; 
    assign layer_0[31] = in[143] ^ in[213]; 
    assign layer_0[32] = ~in[250] | (in[250] & in[132]); 
    assign layer_0[33] = ~(in[189] | in[24]); 
    assign layer_0[34] = in[247] ^ in[203]; 
    assign layer_0[35] = ~(in[89] | in[171]); 
    assign layer_0[36] = ~(in[36] ^ in[178]); 
    assign layer_0[37] = ~in[185] | (in[135] & in[185]); 
    assign layer_0[38] = ~in[76] | (in[76] & in[183]); 
    assign layer_0[39] = in[39] | in[55]; 
    assign layer_0[40] = ~in[11] | (in[92] & in[11]); 
    assign layer_0[41] = ~(in[68] ^ in[80]); 
    assign layer_0[42] = in[93] ^ in[91]; 
    assign layer_0[43] = in[170] ^ in[139]; 
    assign layer_0[44] = in[188] | in[171]; 
    assign layer_0[45] = in[231]; 
    assign layer_0[46] = in[135]; 
    assign layer_0[47] = in[75] & ~in[20]; 
    assign layer_0[48] = in[162] ^ in[180]; 
    assign layer_0[49] = ~(in[90] ^ in[108]); 
    assign layer_0[50] = in[166] & ~in[233]; 
    assign layer_0[51] = in[134] ^ in[185]; 
    assign layer_0[52] = ~(in[195] ^ in[187]); 
    assign layer_0[53] = in[63] ^ in[114]; 
    assign layer_0[54] = in[68] ^ in[71]; 
    assign layer_0[55] = in[251] ^ in[218]; 
    assign layer_0[56] = ~(in[186] ^ in[84]); 
    assign layer_0[57] = ~in[69] | (in[185] & in[69]); 
    assign layer_0[58] = in[58] ^ in[52]; 
    assign layer_0[59] = ~(in[120] | in[76]); 
    assign layer_0[60] = in[131] & ~in[118]; 
    assign layer_0[61] = in[212] ^ in[227]; 
    assign layer_0[62] = in[73]; 
    assign layer_0[63] = in[235]; 
    assign layer_0[64] = ~(in[147] | in[102]); 
    assign layer_0[65] = in[101] | in[70]; 
    assign layer_0[66] = in[243] ^ in[196]; 
    assign layer_0[67] = ~(in[139] & in[136]); 
    assign layer_0[68] = ~(in[242] | in[192]); 
    assign layer_0[69] = ~(in[24] ^ in[72]); 
    assign layer_0[70] = ~(in[119] | in[74]); 
    assign layer_0[71] = ~(in[244] | in[113]); 
    assign layer_0[72] = in[196] ^ in[247]; 
    assign layer_0[73] = ~(in[24] ^ in[27]); 
    assign layer_0[74] = in[56] & ~in[141]; 
    assign layer_0[75] = ~(in[221] ^ in[36]); 
    assign layer_0[76] = in[129] ^ in[131]; 
    assign layer_0[77] = in[132] ^ in[100]; 
    assign layer_0[78] = ~(in[53] ^ in[39]); 
    assign layer_0[79] = in[232] | in[165]; 
    assign layer_0[80] = in[87] ^ in[230]; 
    assign layer_0[81] = ~(in[36] ^ in[68]); 
    assign layer_0[82] = in[103] ^ in[184]; 
    assign layer_0[83] = in[24] ^ in[212]; 
    assign layer_0[84] = in[198] & ~in[136]; 
    assign layer_0[85] = ~(in[116] ^ in[130]); 
    assign layer_0[86] = ~in[123] | (in[123] & in[30]); 
    assign layer_0[87] = in[123] ^ in[137]; 
    assign layer_0[88] = ~in[151] | (in[151] & in[157]); 
    assign layer_0[89] = ~(in[198] | in[212]); 
    assign layer_0[90] = ~in[73]; 
    assign layer_0[91] = in[236] | in[163]; 
    assign layer_0[92] = in[6] ^ in[37]; 
    assign layer_0[93] = in[45] & ~in[41]; 
    assign layer_0[94] = in[91] & in[139]; 
    assign layer_0[95] = in[89] & ~in[211]; 
    assign layer_0[96] = in[9] & ~in[170]; 
    assign layer_0[97] = ~(in[107] | in[89]); 
    assign layer_0[98] = in[219]; 
    assign layer_0[99] = 1'b0; 
    assign layer_0[100] = ~in[153]; 
    assign layer_0[101] = in[41]; 
    assign layer_0[102] = in[93] & ~in[165]; 
    assign layer_0[103] = ~(in[99] ^ in[97]); 
    assign layer_0[104] = ~in[181] | (in[131] & in[181]); 
    assign layer_0[105] = ~(in[67] ^ in[148]); 
    assign layer_0[106] = ~(in[34] | in[91]); 
    assign layer_0[107] = in[247] | in[183]; 
    assign layer_0[108] = in[104] ^ in[87]; 
    assign layer_0[109] = in[7] | in[155]; 
    assign layer_0[110] = in[52] ^ in[155]; 
    assign layer_0[111] = ~(in[119] | in[228]); 
    assign layer_0[112] = ~in[228] | (in[228] & in[23]); 
    assign layer_0[113] = in[23] ^ in[227]; 
    assign layer_0[114] = ~(in[198] ^ in[105]); 
    assign layer_0[115] = ~in[122]; 
    assign layer_0[116] = ~in[90] | (in[78] & in[90]); 
    assign layer_0[117] = ~in[196] | (in[147] & in[196]); 
    assign layer_0[118] = ~(in[241] | in[253]); 
    assign layer_0[119] = ~(in[166] ^ in[132]); 
    assign layer_0[120] = ~(in[91] ^ in[93]); 
    assign layer_0[121] = in[71] | in[40]; 
    assign layer_0[122] = in[24] & ~in[21]; 
    assign layer_0[123] = ~in[252] | (in[252] & in[41]); 
    assign layer_0[124] = in[164] ^ in[153]; 
    assign layer_0[125] = in[21]; 
    assign layer_0[126] = ~in[219]; 
    assign layer_0[127] = in[249] ^ in[203]; 
    assign layer_0[128] = ~(in[120] ^ in[166]); 
    assign layer_0[129] = in[91] & ~in[26]; 
    assign layer_0[130] = ~in[180]; 
    assign layer_0[131] = ~(in[180] | in[143]); 
    assign layer_0[132] = in[163] ^ in[122]; 
    assign layer_0[133] = in[65] | in[90]; 
    assign layer_0[134] = ~in[214] | (in[214] & in[120]); 
    assign layer_0[135] = ~in[245] | (in[172] & in[245]); 
    assign layer_0[136] = in[103] ^ in[116]; 
    assign layer_0[137] = in[221] & ~in[86]; 
    assign layer_0[138] = in[24] & in[71]; 
    assign layer_0[139] = in[110] | in[87]; 
    assign layer_0[140] = ~(in[121] ^ in[89]); 
    assign layer_0[141] = in[170] & ~in[22]; 
    assign layer_0[142] = in[104] ^ in[142]; 
    assign layer_0[143] = ~in[6]; 
    assign layer_0[144] = ~(in[124] ^ in[119]); 
    assign layer_0[145] = in[183] | in[116]; 
    assign layer_0[146] = ~(in[248] ^ in[216]); 
    assign layer_0[147] = ~in[233]; 
    assign layer_0[148] = in[131] | in[199]; 
    assign layer_0[149] = in[125]; 
    assign layer_0[150] = in[249]; 
    assign layer_0[151] = ~(in[50] | in[94]); 
    assign layer_0[152] = in[109] ^ in[111]; 
    assign layer_0[153] = ~(in[88] ^ in[41]); 
    assign layer_0[154] = in[99] | in[70]; 
    assign layer_0[155] = in[119] | in[166]; 
    assign layer_0[156] = in[61] ^ in[27]; 
    assign layer_0[157] = in[211] ^ in[233]; 
    assign layer_0[158] = in[157] | in[155]; 
    assign layer_0[159] = in[83] ^ in[243]; 
    assign layer_0[160] = in[181] & ~in[187]; 
    assign layer_0[161] = in[168] & ~in[52]; 
    assign layer_0[162] = in[81] | in[226]; 
    assign layer_0[163] = in[71] ^ in[24]; 
    assign layer_0[164] = ~(in[215] ^ in[230]); 
    assign layer_0[165] = in[205] ^ in[235]; 
    assign layer_0[166] = in[136] ^ in[117]; 
    assign layer_0[167] = ~(in[170] ^ in[247]); 
    assign layer_0[168] = in[146] & ~in[195]; 
    assign layer_0[169] = in[118] | in[131]; 
    assign layer_0[170] = in[61] | in[66]; 
    assign layer_0[171] = ~(in[28] | in[29]); 
    assign layer_0[172] = in[151] ^ in[119]; 
    assign layer_0[173] = in[200] & ~in[229]; 
    assign layer_0[174] = ~(in[205] | in[164]); 
    assign layer_0[175] = in[197] | in[115]; 
    assign layer_0[176] = ~in[59] | (in[59] & in[84]); 
    assign layer_0[177] = ~(in[68] ^ in[201]); 
    assign layer_0[178] = in[158] | in[198]; 
    assign layer_0[179] = ~(in[180] ^ in[182]); 
    assign layer_0[180] = ~(in[60] | in[155]); 
    assign layer_0[181] = ~(in[39] ^ in[140]); 
    assign layer_0[182] = ~(in[51] ^ in[221]); 
    assign layer_0[183] = ~(in[119] ^ in[90]); 
    assign layer_0[184] = in[178]; 
    assign layer_0[185] = ~(in[117] ^ in[103]); 
    assign layer_0[186] = ~(in[163] | in[99]); 
    assign layer_0[187] = ~(in[35] ^ in[50]); 
    assign layer_0[188] = ~in[12]; 
    assign layer_0[189] = in[9] | in[50]; 
    assign layer_0[190] = ~(in[143] ^ in[157]); 
    assign layer_0[191] = ~in[104] | (in[223] & in[104]); 
    assign layer_0[192] = ~in[99] | (in[99] & in[86]); 
    assign layer_0[193] = ~(in[167] ^ in[243]); 
    assign layer_0[194] = in[166]; 
    assign layer_0[195] = in[140] ^ in[89]; 
    assign layer_0[196] = ~(in[152] | in[120]); 
    assign layer_0[197] = ~(in[88] ^ in[77]); 
    assign layer_0[198] = ~(in[125] | in[46]); 
    assign layer_0[199] = ~in[20]; 
    assign layer_0[200] = ~(in[153] ^ in[82]); 
    assign layer_0[201] = ~(in[182] ^ in[148]); 
    assign layer_0[202] = in[84] & ~in[71]; 
    assign layer_0[203] = in[42] & ~in[138]; 
    assign layer_0[204] = in[120] ^ in[73]; 
    assign layer_0[205] = ~(in[156] | in[180]); 
    assign layer_0[206] = in[215] | in[200]; 
    assign layer_0[207] = in[83] & ~in[177]; 
    assign layer_0[208] = in[177] | in[157]; 
    assign layer_0[209] = ~in[86] | (in[68] & in[86]); 
    assign layer_0[210] = in[235] ^ in[34]; 
    assign layer_0[211] = in[137]; 
    assign layer_0[212] = ~(in[204] | in[76]); 
    assign layer_0[213] = in[114] | in[100]; 
    assign layer_0[214] = ~in[126]; 
    assign layer_0[215] = in[27] | in[194]; 
    assign layer_0[216] = ~(in[98] ^ in[99]); 
    assign layer_0[217] = in[228] | in[40]; 
    assign layer_0[218] = in[238] | in[194]; 
    assign layer_0[219] = ~(in[108] | in[141]); 
    assign layer_0[220] = in[209] ^ in[163]; 
    assign layer_0[221] = ~(in[104] | in[184]); 
    assign layer_0[222] = ~in[120] | (in[120] & in[118]); 
    assign layer_0[223] = ~in[43] | (in[43] & in[106]); 
    assign layer_0[224] = in[167] | in[183]; 
    assign layer_0[225] = ~in[138]; 
    assign layer_0[226] = in[163] & ~in[119]; 
    assign layer_0[227] = ~(in[244] ^ in[165]); 
    assign layer_0[228] = ~in[130] | (in[130] & in[98]); 
    assign layer_0[229] = in[106] & ~in[115]; 
    assign layer_0[230] = ~(in[115] | in[251]); 
    assign layer_0[231] = in[168] & ~in[172]; 
    assign layer_0[232] = ~in[181] | (in[105] & in[181]); 
    assign layer_0[233] = ~(in[203] ^ in[180]); 
    assign layer_0[234] = in[6] | in[27]; 
    assign layer_0[235] = ~(in[119] ^ in[148]); 
    assign layer_0[236] = ~(in[182] ^ in[135]); 
    assign layer_0[237] = ~(in[164] | in[103]); 
    assign layer_0[238] = in[78] | in[54]; 
    assign layer_0[239] = ~(in[134] | in[178]); 
    assign layer_0[240] = in[43] ^ in[73]; 
    assign layer_0[241] = ~(in[248] ^ in[69]); 
    assign layer_0[242] = ~in[21] | (in[243] & in[21]); 
    assign layer_0[243] = ~(in[34] ^ in[66]); 
    assign layer_0[244] = ~(in[69] ^ in[36]); 
    assign layer_0[245] = ~(in[42] | in[213]); 
    assign layer_0[246] = ~(in[131] ^ in[216]); 
    assign layer_0[247] = in[88] ^ in[41]; 
    assign layer_0[248] = ~(in[63] | in[46]); 
    assign layer_0[249] = ~in[248]; 
    assign layer_0[250] = in[137] ^ in[22]; 
    assign layer_0[251] = in[178] | in[27]; 
    assign layer_0[252] = in[197] ^ in[51]; 
    assign layer_0[253] = ~(in[34] | in[243]); 
    assign layer_0[254] = in[117] & in[184]; 
    assign layer_0[255] = in[104] ^ in[166]; 
    assign layer_0[256] = in[121] ^ in[99]; 
    assign layer_0[257] = ~(in[12] ^ in[63]); 
    assign layer_0[258] = ~(in[249] | in[45]); 
    assign layer_0[259] = in[79] | in[87]; 
    assign layer_0[260] = ~(in[168] ^ in[110]); 
    assign layer_0[261] = ~(in[107] & in[106]); 
    assign layer_0[262] = in[148] & ~in[150]; 
    assign layer_0[263] = ~(in[153] ^ in[27]); 
    assign layer_0[264] = in[121] & ~in[179]; 
    assign layer_0[265] = ~(in[83] | in[120]); 
    assign layer_0[266] = ~(in[30] ^ in[79]); 
    assign layer_0[267] = ~(in[115] | in[87]); 
    assign layer_0[268] = in[142] ^ in[24]; 
    assign layer_0[269] = ~(in[179] & in[109]); 
    assign layer_0[270] = in[73] & ~in[151]; 
    assign layer_0[271] = in[181] ^ in[179]; 
    assign layer_0[272] = ~(in[108] ^ in[59]); 
    assign layer_0[273] = ~in[57] | (in[57] & in[131]); 
    assign layer_0[274] = in[214] & ~in[87]; 
    assign layer_0[275] = in[218] ^ in[181]; 
    assign layer_0[276] = ~in[71] | (in[181] & in[71]); 
    assign layer_0[277] = in[60] ^ in[89]; 
    assign layer_0[278] = ~(in[135] | in[54]); 
    assign layer_0[279] = in[85]; 
    assign layer_0[280] = in[252] ^ in[6]; 
    assign layer_0[281] = in[123] ^ in[186]; 
    assign layer_0[282] = in[117] ^ in[130]; 
    assign layer_0[283] = in[83] ^ in[109]; 
    assign layer_0[284] = ~in[54]; 
    assign layer_0[285] = ~(in[110] ^ in[113]); 
    assign layer_0[286] = in[156] | in[92]; 
    assign layer_0[287] = in[232] ^ in[211]; 
    assign layer_0[288] = ~(in[70] ^ in[88]); 
    assign layer_0[289] = in[227] & ~in[40]; 
    assign layer_0[290] = in[176] ^ in[202]; 
    assign layer_0[291] = ~(in[196] ^ in[130]); 
    assign layer_0[292] = ~(in[90] | in[58]); 
    assign layer_0[293] = in[59] | in[75]; 
    assign layer_0[294] = ~(in[89] | in[110]); 
    assign layer_0[295] = in[73] & ~in[21]; 
    assign layer_0[296] = in[91] ^ in[78]; 
    assign layer_0[297] = in[219]; 
    assign layer_0[298] = ~(in[159] | in[186]); 
    assign layer_0[299] = in[102]; 
    assign layer_0[300] = in[7] | in[214]; 
    assign layer_0[301] = ~(in[250] ^ in[202]); 
    assign layer_0[302] = in[90] | in[70]; 
    assign layer_0[303] = ~(in[170] ^ in[167]); 
    assign layer_0[304] = in[245] & ~in[25]; 
    assign layer_0[305] = ~(in[41] ^ in[88]); 
    assign layer_0[306] = in[152] ^ in[183]; 
    assign layer_0[307] = ~(in[231] ^ in[216]); 
    assign layer_0[308] = in[212] | in[58]; 
    assign layer_0[309] = in[158] & ~in[87]; 
    assign layer_0[310] = ~in[85]; 
    assign layer_0[311] = ~in[60]; 
    assign layer_0[312] = ~in[40]; 
    assign layer_0[313] = ~(in[136] ^ in[249]); 
    assign layer_0[314] = in[9]; 
    assign layer_0[315] = ~in[182] | (in[110] & in[182]); 
    assign layer_0[316] = ~(in[164] | in[181]); 
    assign layer_0[317] = ~(in[165] ^ in[202]); 
    assign layer_0[318] = in[149] ^ in[151]; 
    assign layer_0[319] = ~(in[249] ^ in[100]); 
    assign layer_0[320] = in[82] ^ in[105]; 
    assign layer_0[321] = in[57] & ~in[219]; 
    assign layer_0[322] = in[197] ^ in[245]; 
    assign layer_0[323] = ~(in[79] ^ in[47]); 
    assign layer_0[324] = ~(in[126] | in[127]); 
    assign layer_0[325] = in[11] ^ in[206]; 
    assign layer_0[326] = in[217] ^ in[211]; 
    assign layer_0[327] = in[186] | in[53]; 
    assign layer_0[328] = ~(in[214] & in[134]); 
    assign layer_0[329] = ~(in[230] | in[195]); 
    assign layer_0[330] = in[249] ^ in[236]; 
    assign layer_0[331] = in[102] | in[79]; 
    assign layer_0[332] = in[137] ^ in[154]; 
    assign layer_0[333] = ~(in[55] ^ in[53]); 
    assign layer_0[334] = ~(in[55] ^ in[39]); 
    assign layer_0[335] = ~(in[125] ^ in[134]); 
    assign layer_0[336] = ~in[135]; 
    assign layer_0[337] = in[26] | in[108]; 
    assign layer_0[338] = ~(in[52] ^ in[106]); 
    assign layer_0[339] = ~(in[60] | in[52]); 
    assign layer_0[340] = ~(in[54] ^ in[7]); 
    assign layer_0[341] = in[197] | in[94]; 
    assign layer_0[342] = ~(in[107] ^ in[139]); 
    assign layer_0[343] = ~in[171] | (in[171] & in[104]); 
    assign layer_0[344] = ~(in[155] | in[12]); 
    assign layer_0[345] = in[235] ^ in[89]; 
    assign layer_0[346] = in[76] | in[211]; 
    assign layer_0[347] = ~(in[60] ^ in[72]); 
    assign layer_0[348] = ~(in[117] | in[102]); 
    assign layer_0[349] = in[119] & ~in[60]; 
    assign layer_0[350] = ~(in[223] ^ in[253]); 
    assign layer_0[351] = ~in[130] | (in[135] & in[130]); 
    assign layer_0[352] = in[198] ^ in[216]; 
    assign layer_0[353] = in[142]; 
    assign layer_0[354] = in[6] | in[50]; 
    assign layer_0[355] = in[199] & ~in[245]; 
    assign layer_0[356] = in[135] | in[150]; 
    assign layer_0[357] = ~(in[185] ^ in[188]); 
    assign layer_0[358] = ~(in[146] ^ in[148]); 
    assign layer_0[359] = in[228] & ~in[30]; 
    assign layer_0[360] = ~(in[172] | in[198]); 
    assign layer_0[361] = ~(in[184] ^ in[230]); 
    assign layer_0[362] = in[156] & in[72]; 
    assign layer_0[363] = ~(in[87] ^ in[72]); 
    assign layer_0[364] = in[84] ^ in[181]; 
    assign layer_0[365] = ~(in[141] ^ in[19]); 
    assign layer_0[366] = in[135]; 
    assign layer_0[367] = in[219] ^ in[173]; 
    assign layer_0[368] = in[163] ^ in[184]; 
    assign layer_0[369] = ~in[134]; 
    assign layer_0[370] = ~in[51]; 
    assign layer_0[371] = in[88] ^ in[119]; 
    assign layer_0[372] = in[105] ^ in[169]; 
    assign layer_0[373] = ~in[113]; 
    assign layer_0[374] = ~in[165]; 
    assign layer_0[375] = in[129] ^ in[137]; 
    assign layer_0[376] = ~(in[214] ^ in[229]); 
    assign layer_0[377] = ~(in[28] | in[92]); 
    assign layer_0[378] = ~(in[125] & in[114]); 
    assign layer_0[379] = ~in[140]; 
    assign layer_0[380] = in[75] | in[76]; 
    assign layer_0[381] = ~(in[78] ^ in[206]); 
    assign layer_0[382] = in[39] | in[59]; 
    assign layer_0[383] = ~(in[111] ^ in[109]); 
    assign layer_0[384] = ~(in[197] ^ in[85]); 
    assign layer_0[385] = ~in[104] | (in[104] & in[135]); 
    assign layer_0[386] = in[90] ^ in[122]; 
    assign layer_0[387] = in[68] & ~in[211]; 
    assign layer_0[388] = ~in[135] | (in[135] & in[139]); 
    assign layer_0[389] = ~(in[242] | in[22]); 
    assign layer_0[390] = ~(in[101] | in[92]); 
    assign layer_0[391] = ~(in[225] ^ in[246]); 
    assign layer_0[392] = in[181] ^ in[85]; 
    assign layer_0[393] = in[126] ^ in[125]; 
    assign layer_0[394] = ~(in[172] | in[179]); 
    assign layer_0[395] = ~(in[177] | in[26]); 
    assign layer_0[396] = ~(in[110] ^ in[108]); 
    assign layer_0[397] = ~(in[180] | in[217]); 
    assign layer_0[398] = ~in[71] | (in[71] & in[227]); 
    assign layer_0[399] = ~(in[135] | in[251]); 
    assign layer_0[400] = in[58] & ~in[200]; 
    assign layer_0[401] = ~(in[209] ^ in[143]); 
    assign layer_0[402] = in[187] ^ in[232]; 
    assign layer_0[403] = ~in[198] | (in[198] & in[220]); 
    assign layer_0[404] = ~(in[131] ^ in[133]); 
    assign layer_0[405] = ~in[75] | (in[220] & in[75]); 
    assign layer_0[406] = in[149] ^ in[117]; 
    assign layer_0[407] = in[91] ^ in[56]; 
    assign layer_0[408] = in[110] & ~in[231]; 
    assign layer_0[409] = in[221] ^ in[249]; 
    assign layer_0[410] = in[57] & ~in[157]; 
    assign layer_0[411] = ~(in[67] ^ in[117]); 
    assign layer_0[412] = in[23] | in[93]; 
    assign layer_0[413] = ~(in[77] ^ in[78]); 
    assign layer_0[414] = in[73] ^ in[88]; 
    assign layer_0[415] = ~(in[21] ^ in[85]); 
    assign layer_0[416] = in[230] & ~in[178]; 
    assign layer_0[417] = in[134] & ~in[13]; 
    assign layer_0[418] = ~(in[234] | in[196]); 
    assign layer_0[419] = in[197]; 
    assign layer_0[420] = in[146] ^ in[163]; 
    assign layer_0[421] = ~(in[46] ^ in[236]); 
    assign layer_0[422] = ~(in[233] | in[211]); 
    assign layer_0[423] = ~(in[155] | in[177]); 
    assign layer_0[424] = ~(in[97] ^ in[77]); 
    assign layer_0[425] = ~in[143]; 
    assign layer_0[426] = ~in[89] | (in[89] & in[27]); 
    assign layer_0[427] = ~(in[167] ^ in[99]); 
    assign layer_0[428] = ~(in[182] ^ in[164]); 
    assign layer_0[429] = ~(in[123] ^ in[140]); 
    assign layer_0[430] = in[46] ^ in[29]; 
    assign layer_0[431] = in[249]; 
    assign layer_0[432] = in[130]; 
    assign layer_0[433] = ~(in[132] | in[10]); 
    assign layer_0[434] = in[136] | in[197]; 
    assign layer_0[435] = ~(in[206] ^ in[236]); 
    assign layer_0[436] = ~in[30] | (in[30] & in[92]); 
    assign layer_0[437] = in[78] | in[231]; 
    assign layer_0[438] = in[106] & ~in[61]; 
    assign layer_0[439] = in[85] | in[93]; 
    assign layer_0[440] = ~in[78]; 
    assign layer_0[441] = in[166] | in[24]; 
    assign layer_0[442] = ~(in[51] ^ in[229]); 
    assign layer_0[443] = ~(in[142] | in[132]); 
    assign layer_0[444] = ~in[103] | (in[103] & in[84]); 
    assign layer_0[445] = ~(in[109] | in[136]); 
    assign layer_0[446] = in[153] ^ in[122]; 
    assign layer_0[447] = ~(in[151] ^ in[182]); 
    assign layer_0[448] = ~in[75]; 
    assign layer_0[449] = ~(in[148] ^ in[134]); 
    assign layer_0[450] = in[249] ^ in[215]; 
    assign layer_0[451] = in[57] & ~in[155]; 
    assign layer_0[452] = ~(in[88] | in[9]); 
    assign layer_0[453] = in[25] ^ in[28]; 
    assign layer_0[454] = ~(in[51] ^ in[11]); 
    assign layer_0[455] = ~(in[53] | in[38]); 
    assign layer_0[456] = ~(in[52] ^ in[83]); 
    assign layer_0[457] = in[150] ^ in[98]; 
    assign layer_0[458] = ~in[143]; 
    assign layer_0[459] = ~in[122]; 
    assign layer_0[460] = in[115] & ~in[188]; 
    assign layer_0[461] = in[57] ^ in[41]; 
    assign layer_0[462] = ~(in[140] ^ in[141]); 
    assign layer_0[463] = ~(in[204] ^ in[236]); 
    assign layer_0[464] = in[178] | in[231]; 
    assign layer_0[465] = in[133] | in[116]; 
    assign layer_0[466] = ~(in[231] | in[94]); 
    assign layer_0[467] = in[135] ^ in[101]; 
    assign layer_0[468] = in[52] | in[91]; 
    assign layer_0[469] = in[197] ^ in[228]; 
    assign layer_0[470] = in[92] | in[105]; 
    assign layer_0[471] = ~(in[98] ^ in[87]); 
    assign layer_0[472] = in[56] | in[72]; 
    assign layer_0[473] = in[235]; 
    assign layer_0[474] = ~in[51] | (in[35] & in[51]); 
    assign layer_0[475] = in[119] ^ in[133]; 
    assign layer_0[476] = ~in[153] | (in[153] & in[59]); 
    assign layer_0[477] = ~(in[122] ^ in[156]); 
    assign layer_0[478] = in[72] | in[40]; 
    assign layer_0[479] = in[88] ^ in[132]; 
    assign layer_0[480] = in[106] ^ in[108]; 
    assign layer_0[481] = in[99] | in[150]; 
    assign layer_0[482] = in[100] ^ in[105]; 
    assign layer_0[483] = ~in[56] | (in[8] & in[56]); 
    assign layer_0[484] = in[152] | in[183]; 
    assign layer_0[485] = in[235]; 
    assign layer_0[486] = in[125] | in[155]; 
    assign layer_0[487] = ~in[167]; 
    assign layer_0[488] = ~(in[182] ^ in[185]); 
    assign layer_0[489] = in[133]; 
    assign layer_0[490] = in[9] ^ in[12]; 
    assign layer_0[491] = ~(in[213] ^ in[244]); 
    assign layer_0[492] = in[164] ^ in[182]; 
    assign layer_0[493] = ~(in[58] | in[71]); 
    assign layer_0[494] = ~(in[20] | in[179]); 
    assign layer_0[495] = in[217] ^ in[249]; 
    assign layer_0[496] = ~(in[155] | in[99]); 
    assign layer_0[497] = in[116]; 
    assign layer_0[498] = in[45] ^ in[76]; 
    assign layer_0[499] = ~(in[50] ^ in[248]); 
    assign layer_0[500] = ~(in[109] | in[39]); 
    assign layer_0[501] = in[181] & ~in[107]; 
    assign layer_0[502] = in[117] | in[34]; 
    assign layer_0[503] = in[248]; 
    assign layer_0[504] = in[248] & ~in[214]; 
    assign layer_0[505] = in[7] ^ in[214]; 
    assign layer_0[506] = in[135] ^ in[166]; 
    assign layer_0[507] = ~(in[76] ^ in[120]); 
    assign layer_0[508] = in[74] & ~in[56]; 
    assign layer_0[509] = in[165] | in[178]; 
    assign layer_0[510] = in[97] | in[247]; 
    assign layer_0[511] = in[87] ^ in[100]; 
    assign layer_0[512] = ~(in[98] ^ in[183]); 
    assign layer_0[513] = in[148] ^ in[130]; 
    assign layer_0[514] = ~(in[9] ^ in[148]); 
    assign layer_0[515] = ~(in[125] | in[102]); 
    assign layer_0[516] = ~(in[108] ^ in[90]); 
    assign layer_0[517] = in[121] ^ in[250]; 
    assign layer_0[518] = in[99] ^ in[117]; 
    assign layer_0[519] = in[231] | in[231]; 
    assign layer_0[520] = ~(in[50] | in[20]); 
    assign layer_0[521] = in[170] & ~in[213]; 
    assign layer_0[522] = in[30]; 
    assign layer_0[523] = ~(in[218] ^ in[183]); 
    assign layer_0[524] = ~in[72] | (in[72] & in[47]); 
    assign layer_0[525] = ~(in[56] ^ in[25]); 
    assign layer_0[526] = ~(in[181] ^ in[85]); 
    assign layer_0[527] = ~(in[170] ^ in[227]); 
    assign layer_0[528] = ~(in[180] | in[195]); 
    assign layer_0[529] = ~(in[214] ^ in[22]); 
    assign layer_0[530] = in[185] ^ in[235]; 
    assign layer_0[531] = in[75] ^ in[106]; 
    assign layer_0[532] = ~in[169]; 
    assign layer_0[533] = ~(in[235] | in[212]); 
    assign layer_0[534] = ~(in[228] ^ in[198]); 
    assign layer_0[535] = ~(in[108] | in[110]); 
    assign layer_0[536] = ~in[189]; 
    assign layer_0[537] = in[185] ^ in[150]; 
    assign layer_0[538] = in[162] ^ in[104]; 
    assign layer_0[539] = ~(in[99] ^ in[101]); 
    assign layer_0[540] = ~(in[140] | in[122]); 
    assign layer_0[541] = in[217] ^ in[249]; 
    assign layer_0[542] = ~(in[236] | in[201]); 
    assign layer_0[543] = ~(in[251] | in[51]); 
    assign layer_0[544] = in[46] | in[235]; 
    assign layer_0[545] = in[20] | in[186]; 
    assign layer_0[546] = ~in[86]; 
    assign layer_0[547] = ~in[41]; 
    assign layer_0[548] = ~(in[120] | in[245]); 
    assign layer_0[549] = in[151] | in[93]; 
    assign layer_0[550] = ~(in[213] ^ in[245]); 
    assign layer_0[551] = in[53] ^ in[92]; 
    assign layer_0[552] = ~(in[85] ^ in[36]); 
    assign layer_0[553] = in[236]; 
    assign layer_0[554] = in[86]; 
    assign layer_0[555] = ~in[105]; 
    assign layer_0[556] = ~(in[140] ^ in[126]); 
    assign layer_0[557] = in[188] | in[149]; 
    assign layer_0[558] = in[103] ^ in[116]; 
    assign layer_0[559] = in[149] ^ in[183]; 
    assign layer_0[560] = in[246] | in[214]; 
    assign layer_0[561] = in[51] | in[194]; 
    assign layer_0[562] = in[210] | in[37]; 
    assign layer_0[563] = ~(in[71] ^ in[170]); 
    assign layer_0[564] = in[143] ^ in[27]; 
    assign layer_0[565] = ~(in[91] ^ in[102]); 
    assign layer_0[566] = in[168] & ~in[177]; 
    assign layer_0[567] = in[93]; 
    assign layer_0[568] = ~in[56] | (in[101] & in[56]); 
    assign layer_0[569] = in[141] ^ in[139]; 
    assign layer_0[570] = in[59] ^ in[55]; 
    assign layer_0[571] = ~in[180]; 
    assign layer_0[572] = ~(in[120] | in[88]); 
    assign layer_0[573] = in[120] & ~in[172]; 
    assign layer_0[574] = in[133] & ~in[107]; 
    assign layer_0[575] = ~in[148] | (in[98] & in[148]); 
    assign layer_0[576] = in[244] | in[231]; 
    assign layer_0[577] = in[242] | in[8]; 
    assign layer_0[578] = in[199] ^ in[186]; 
    assign layer_0[579] = ~(in[165] ^ in[167]); 
    assign layer_0[580] = ~(in[155] | in[86]); 
    assign layer_0[581] = in[103] ^ in[117]; 
    assign layer_0[582] = ~(in[202] ^ in[51]); 
    assign layer_0[583] = ~(in[121] ^ in[153]); 
    assign layer_0[584] = in[217]; 
    assign layer_0[585] = in[59] & ~in[106]; 
    assign layer_0[586] = in[142] | in[169]; 
    assign layer_0[587] = ~in[179]; 
    assign layer_0[588] = in[168] | in[137]; 
    assign layer_0[589] = in[141]; 
    assign layer_0[590] = ~(in[67] ^ in[35]); 
    assign layer_0[591] = ~(in[250] | in[167]); 
    assign layer_0[592] = in[36] ^ in[104]; 
    assign layer_0[593] = ~(in[38] | in[187]); 
    assign layer_0[594] = in[148] ^ in[119]; 
    assign layer_0[595] = ~(in[22] ^ in[53]); 
    assign layer_0[596] = ~in[182]; 
    assign layer_0[597] = in[59] ^ in[235]; 
    assign layer_0[598] = in[223] | in[8]; 
    assign layer_0[599] = in[154] & ~in[221]; 
    assign layer_0[600] = ~(in[91] | in[183]); 
    assign layer_0[601] = ~(in[175] | in[162]); 
    assign layer_0[602] = ~(in[106] | in[138]); 
    assign layer_0[603] = ~in[117] | (in[117] & in[151]); 
    assign layer_0[604] = ~(in[95] | in[11]); 
    assign layer_0[605] = ~in[58] | (in[121] & in[58]); 
    assign layer_0[606] = ~(in[35] | in[132]); 
    assign layer_0[607] = in[106] ^ in[108]; 
    assign layer_0[608] = in[115] ^ in[116]; 
    assign layer_0[609] = ~in[44] | (in[70] & in[44]); 
    assign layer_0[610] = ~(in[105] ^ in[43]); 
    assign layer_0[611] = ~(in[109] & in[110]); 
    assign layer_0[612] = in[159] | in[183]; 
    assign layer_0[613] = ~(in[100] ^ in[102]); 
    assign layer_0[614] = ~(in[68] | in[120]); 
    assign layer_0[615] = ~in[86] | (in[22] & in[86]); 
    assign layer_0[616] = ~(in[163] ^ in[109]); 
    assign layer_0[617] = ~in[151] | (in[151] & in[86]); 
    assign layer_0[618] = ~(in[211] | in[104]); 
    assign layer_0[619] = ~in[248] | (in[248] & in[169]); 
    assign layer_0[620] = in[67] | in[184]; 
    assign layer_0[621] = in[150]; 
    assign layer_0[622] = ~(in[42] ^ in[86]); 
    assign layer_0[623] = ~(in[249] ^ in[236]); 
    assign layer_0[624] = in[133] | in[151]; 
    assign layer_0[625] = in[134] ^ in[235]; 
    assign layer_0[626] = ~(in[24] ^ in[196]); 
    assign layer_0[627] = 1'b0; 
    assign layer_0[628] = in[151] ^ in[122]; 
    assign layer_0[629] = ~(in[245] | in[247]); 
    assign layer_0[630] = ~(in[6] ^ in[188]); 
    assign layer_0[631] = in[10] | in[12]; 
    assign layer_0[632] = ~in[153] | (in[179] & in[153]); 
    assign layer_0[633] = in[41] ^ in[71]; 
    assign layer_0[634] = ~in[40] | (in[10] & in[40]); 
    assign layer_0[635] = in[69] | in[91]; 
    assign layer_0[636] = in[26] ^ in[59]; 
    assign layer_0[637] = in[165] ^ in[213]; 
    assign layer_0[638] = ~(in[105] | in[162]); 
    assign layer_0[639] = in[38] ^ in[247]; 
    assign layer_0[640] = ~in[198] | (in[198] & in[210]); 
    assign layer_0[641] = ~in[120] | (in[162] & in[120]); 
    assign layer_0[642] = in[219] | in[204]; 
    assign layer_0[643] = ~(in[143] | in[195]); 
    assign layer_0[644] = in[91] ^ in[77]; 
    assign layer_0[645] = ~(in[89] ^ in[104]); 
    assign layer_0[646] = in[140] ^ in[87]; 
    assign layer_0[647] = in[57] & ~in[213]; 
    assign layer_0[648] = in[102] ^ in[129]; 
    assign layer_0[649] = in[129] ^ in[101]; 
    assign layer_0[650] = ~(in[136] ^ in[70]); 
    assign layer_0[651] = ~in[57] | (in[54] & in[57]); 
    assign layer_0[652] = in[30] ^ in[215]; 
    assign layer_0[653] = ~in[165]; 
    assign layer_0[654] = ~in[250] | (in[250] & in[188]); 
    assign layer_0[655] = in[170]; 
    assign layer_0[656] = in[162] ^ in[165]; 
    assign layer_0[657] = in[159] ^ in[213]; 
    assign layer_0[658] = ~in[244]; 
    assign layer_0[659] = in[95] | in[83]; 
    assign layer_0[660] = ~in[79]; 
    assign layer_0[661] = ~in[54] | (in[140] & in[54]); 
    assign layer_0[662] = ~(in[221] ^ in[154]); 
    assign layer_0[663] = ~in[140] | (in[140] & in[60]); 
    assign layer_0[664] = in[221] ^ in[69]; 
    assign layer_0[665] = ~in[115] | (in[195] & in[115]); 
    assign layer_0[666] = in[168] ^ in[248]; 
    assign layer_0[667] = in[233] ^ in[231]; 
    assign layer_0[668] = ~(in[26] | in[29]); 
    assign layer_0[669] = in[153] & ~in[8]; 
    assign layer_0[670] = in[138] ^ in[187]; 
    assign layer_0[671] = in[115] & ~in[120]; 
    assign layer_0[672] = in[154] & ~in[196]; 
    assign layer_0[673] = ~(in[154] ^ in[24]); 
    assign layer_0[674] = ~(in[198] ^ in[245]); 
    assign layer_0[675] = in[143] ^ in[196]; 
    assign layer_0[676] = in[134] ^ in[103]; 
    assign layer_0[677] = ~(in[187] | in[225]); 
    assign layer_0[678] = ~(in[75] ^ in[106]); 
    assign layer_0[679] = ~(in[42] ^ in[123]); 
    assign layer_0[680] = in[9] & ~in[232]; 
    assign layer_0[681] = in[62] ^ in[44]; 
    assign layer_0[682] = ~in[157] | (in[157] & in[86]); 
    assign layer_0[683] = in[244] | in[24]; 
    assign layer_0[684] = in[106] | in[67]; 
    assign layer_0[685] = ~in[149]; 
    assign layer_0[686] = ~(in[183] | in[180]); 
    assign layer_0[687] = in[84] | in[108]; 
    assign layer_0[688] = in[167]; 
    assign layer_0[689] = ~(in[152] ^ in[199]); 
    assign layer_0[690] = ~(in[232] ^ in[183]); 
    assign layer_0[691] = in[163] | in[157]; 
    assign layer_0[692] = in[28]; 
    assign layer_0[693] = in[102]; 
    assign layer_0[694] = in[170] ^ in[250]; 
    assign layer_0[695] = ~(in[25] ^ in[44]); 
    assign layer_0[696] = ~(in[252] ^ in[149]); 
    assign layer_0[697] = ~(in[30] ^ in[79]); 
    assign layer_0[698] = ~(in[97] ^ in[99]); 
    assign layer_0[699] = ~(in[202] ^ in[234]); 
    assign layer_0[700] = ~(in[250] ^ in[70]); 
    assign layer_0[701] = in[154] & ~in[77]; 
    assign layer_0[702] = ~(in[95] | in[45]); 
    assign layer_0[703] = ~(in[195] | in[198]); 
    assign layer_0[704] = in[73] ^ in[75]; 
    assign layer_0[705] = ~(in[109] | in[124]); 
    assign layer_0[706] = in[86] & ~in[41]; 
    assign layer_0[707] = ~(in[225] | in[105]); 
    assign layer_0[708] = ~(in[132] | in[143]); 
    assign layer_0[709] = ~in[36] | (in[103] & in[36]); 
    assign layer_0[710] = in[156] | in[230]; 
    assign layer_0[711] = in[165] | in[167]; 
    assign layer_0[712] = in[204] ^ in[140]; 
    assign layer_0[713] = in[19] ^ in[101]; 
    assign layer_0[714] = ~(in[77] ^ in[90]); 
    assign layer_0[715] = ~(in[130] ^ in[57]); 
    assign layer_0[716] = in[165] ^ in[69]; 
    assign layer_0[717] = ~(in[167] | in[237]); 
    assign layer_0[718] = ~(in[119] ^ in[232]); 
    assign layer_0[719] = ~(in[93] ^ in[73]); 
    assign layer_0[720] = in[210] | in[61]; 
    assign layer_0[721] = ~in[165] | (in[165] & in[169]); 
    assign layer_0[722] = in[136] ^ in[167]; 
    assign layer_0[723] = in[184] & ~in[54]; 
    assign layer_0[724] = ~(in[85] ^ in[39]); 
    assign layer_0[725] = ~in[89] | (in[89] & in[10]); 
    assign layer_0[726] = ~(in[164] | in[181]); 
    assign layer_0[727] = ~(in[248] | in[136]); 
    assign layer_0[728] = in[95] | in[79]; 
    assign layer_0[729] = in[173] ^ in[205]; 
    assign layer_0[730] = in[119] & ~in[186]; 
    assign layer_0[731] = in[121] & in[122]; 
    assign layer_0[732] = ~(in[183] ^ in[77]); 
    assign layer_0[733] = in[98] | in[101]; 
    assign layer_0[734] = ~(in[98] | in[38]); 
    assign layer_0[735] = ~(in[156] | in[100]); 
    assign layer_0[736] = in[110] ^ in[92]; 
    assign layer_0[737] = in[25] ^ in[93]; 
    assign layer_0[738] = in[68] ^ in[86]; 
    assign layer_0[739] = ~(in[231] | in[228]); 
    assign layer_0[740] = in[175] ^ in[218]; 
    assign layer_0[741] = in[31] | in[76]; 
    assign layer_0[742] = ~in[181]; 
    assign layer_0[743] = in[242] ^ in[248]; 
    assign layer_0[744] = ~(in[82] | in[158]); 
    assign layer_0[745] = ~in[234]; 
    assign layer_0[746] = in[97] ^ in[103]; 
    assign layer_0[747] = ~(in[117] ^ in[131]); 
    assign layer_0[748] = in[153] & ~in[237]; 
    assign layer_0[749] = ~(in[237] ^ in[82]); 
    assign layer_0[750] = in[137] & ~in[232]; 
    assign layer_0[751] = ~in[193]; 
    assign layer_0[752] = in[57] & ~in[37]; 
    assign layer_0[753] = ~in[181]; 
    assign layer_0[754] = ~(in[135] ^ in[102]); 
    assign layer_0[755] = ~(in[124] | in[91]); 
    assign layer_0[756] = in[138] & ~in[204]; 
    assign layer_0[757] = ~(in[104] ^ in[74]); 
    assign layer_0[758] = in[193] | in[47]; 
    assign layer_0[759] = in[185] | in[146]; 
    assign layer_0[760] = ~(in[56] | in[72]); 
    assign layer_0[761] = ~(in[28] ^ in[194]); 
    assign layer_0[762] = ~(in[107] ^ in[124]); 
    assign layer_0[763] = in[186] & ~in[235]; 
    assign layer_0[764] = in[23] ^ in[186]; 
    assign layer_0[765] = ~in[70] | (in[70] & in[68]); 
    assign layer_0[766] = in[137] & ~in[214]; 
    assign layer_0[767] = in[121] & ~in[219]; 
    assign layer_0[768] = ~in[57] | (in[152] & in[57]); 
    assign layer_0[769] = in[104] ^ in[74]; 
    assign layer_0[770] = in[154] & ~in[59]; 
    assign layer_0[771] = ~(in[195] | in[135]); 
    assign layer_0[772] = in[177] | in[222]; 
    assign layer_0[773] = in[167] ^ in[108]; 
    assign layer_0[774] = in[180] ^ in[150]; 
    assign layer_0[775] = in[165] ^ in[101]; 
    assign layer_0[776] = ~in[146] | (in[146] & in[120]); 
    assign layer_0[777] = in[219] | in[204]; 
    assign layer_0[778] = ~(in[38] ^ in[66]); 
    assign layer_0[779] = ~(in[116] | in[118]); 
    assign layer_0[780] = in[105] | in[106]; 
    assign layer_0[781] = in[110] ^ in[109]; 
    assign layer_0[782] = in[177] ^ in[190]; 
    assign layer_0[783] = in[20] ^ in[90]; 
    assign layer_0[784] = in[196] ^ in[165]; 
    assign layer_0[785] = in[217] & ~in[249]; 
    assign layer_0[786] = ~(in[163] | in[27]); 
    assign layer_0[787] = in[46] ^ in[234]; 
    assign layer_0[788] = in[90] | in[69]; 
    assign layer_0[789] = in[52] ^ in[58]; 
    assign layer_0[790] = in[170]; 
    assign layer_0[791] = ~(in[197] ^ in[85]); 
    assign layer_0[792] = in[61] | in[146]; 
    assign layer_0[793] = ~(in[108] | in[93]); 
    assign layer_0[794] = ~(in[127] ^ in[43]); 
    assign layer_0[795] = in[68] ^ in[105]; 
    assign layer_0[796] = in[165]; 
    assign layer_0[797] = ~(in[69] ^ in[170]); 
    assign layer_0[798] = ~(in[245] | in[250]); 
    assign layer_0[799] = in[179] | in[180]; 
    assign layer_0[800] = in[182]; 
    assign layer_0[801] = in[155] | in[198]; 
    assign layer_0[802] = in[55] | in[45]; 
    assign layer_0[803] = ~in[19]; 
    assign layer_0[804] = ~(in[216] ^ in[195]); 
    assign layer_0[805] = in[189] | in[245]; 
    assign layer_0[806] = ~(in[161] | in[223]); 
    assign layer_0[807] = ~(in[31] ^ in[74]); 
    assign layer_0[808] = in[196] ^ in[204]; 
    assign layer_0[809] = in[102] ^ in[84]; 
    assign layer_0[810] = in[91] | in[164]; 
    assign layer_0[811] = ~in[84] | (in[84] & in[137]); 
    assign layer_0[812] = ~in[116] | (in[116] & in[183]); 
    assign layer_0[813] = in[150] | in[180]; 
    assign layer_0[814] = ~(in[163] | in[215]); 
    assign layer_0[815] = ~(in[131] ^ in[167]); 
    assign layer_0[816] = in[186] & ~in[197]; 
    assign layer_0[817] = in[74] & ~in[125]; 
    assign layer_0[818] = in[8]; 
    assign layer_0[819] = ~(in[195] | in[38]); 
    assign layer_0[820] = ~(in[91] ^ in[93]); 
    assign layer_0[821] = ~(in[195] | in[4]); 
    assign layer_0[822] = in[122] & ~in[170]; 
    assign layer_0[823] = in[91] ^ in[109]; 
    assign layer_0[824] = ~(in[91] ^ in[93]); 
    assign layer_0[825] = ~(in[7] ^ in[219]); 
    assign layer_0[826] = in[113] | in[114]; 
    assign layer_0[827] = ~(in[34] ^ in[104]); 
    assign layer_0[828] = in[118] & ~in[24]; 
    assign layer_0[829] = ~in[89] | (in[89] & in[135]); 
    assign layer_0[830] = in[58] ^ in[29]; 
    assign layer_0[831] = ~in[120] | (in[120] & in[168]); 
    assign layer_0[832] = in[72] | in[93]; 
    assign layer_0[833] = in[71] ^ in[212]; 
    assign layer_0[834] = in[9] ^ in[63]; 
    assign layer_0[835] = ~(in[148] ^ in[183]); 
    assign layer_0[836] = in[207] | in[26]; 
    assign layer_0[837] = ~in[183] | (in[250] & in[183]); 
    assign layer_0[838] = ~(in[130] ^ in[180]); 
    assign layer_0[839] = ~in[103] | (in[170] & in[103]); 
    assign layer_0[840] = in[253] | in[202]; 
    assign layer_0[841] = in[115]; 
    assign layer_0[842] = ~(in[118] ^ in[113]); 
    assign layer_0[843] = ~(in[27] ^ in[24]); 
    assign layer_0[844] = ~(in[199] ^ in[89]); 
    assign layer_0[845] = in[213] & ~in[156]; 
    assign layer_0[846] = in[105] & in[118]; 
    assign layer_0[847] = ~(in[195] ^ in[250]); 
    assign layer_0[848] = ~in[41]; 
    assign layer_0[849] = in[70] ^ in[22]; 
    assign layer_0[850] = ~(in[86] ^ in[72]); 
    assign layer_0[851] = in[228] | in[199]; 
    assign layer_0[852] = ~(in[6] | in[120]); 
    assign layer_0[853] = ~(in[103] ^ in[56]); 
    assign layer_0[854] = ~(in[105] ^ in[26]); 
    assign layer_0[855] = ~(in[201] | in[164]); 
    assign layer_0[856] = in[230]; 
    assign layer_0[857] = in[60] | in[86]; 
    assign layer_0[858] = in[87] ^ in[24]; 
    assign layer_0[859] = ~(in[209] | in[109]); 
    assign layer_0[860] = ~(in[41] | in[56]); 
    assign layer_0[861] = ~in[86]; 
    assign layer_0[862] = ~(in[19] ^ in[102]); 
    assign layer_0[863] = ~(in[221] ^ in[212]); 
    assign layer_0[864] = ~(in[75] ^ in[42]); 
    assign layer_0[865] = ~(in[155] | in[162]); 
    assign layer_0[866] = in[61] | in[40]; 
    assign layer_0[867] = in[94] & ~in[243]; 
    assign layer_0[868] = in[85] | in[196]; 
    assign layer_0[869] = in[228] ^ in[56]; 
    assign layer_0[870] = ~(in[118] ^ in[173]); 
    assign layer_0[871] = ~in[126]; 
    assign layer_0[872] = in[194] | in[179]; 
    assign layer_0[873] = ~(in[70] ^ in[201]); 
    assign layer_0[874] = in[41] | in[9]; 
    assign layer_0[875] = ~(in[103] ^ in[70]); 
    assign layer_0[876] = in[73] | in[94]; 
    assign layer_0[877] = ~in[213] | (in[213] & in[137]); 
    assign layer_0[878] = ~in[76]; 
    assign layer_0[879] = in[86]; 
    assign layer_0[880] = ~(in[219] | in[132]); 
    assign layer_0[881] = ~(in[158] ^ in[108]); 
    assign layer_0[882] = in[164] ^ in[135]; 
    assign layer_0[883] = ~(in[104] | in[180]); 
    assign layer_0[884] = ~(in[44] ^ in[42]); 
    assign layer_0[885] = ~(in[132] & in[132]); 
    assign layer_0[886] = ~(in[198] ^ in[228]); 
    assign layer_0[887] = ~in[168] | (in[165] & in[168]); 
    assign layer_0[888] = ~(in[148] & in[54]); 
    assign layer_0[889] = in[148] ^ in[150]; 
    assign layer_0[890] = in[39] & ~in[227]; 
    assign layer_0[891] = in[40] ^ in[71]; 
    assign layer_0[892] = ~(in[193] | in[242]); 
    assign layer_0[893] = ~(in[147] | in[154]); 
    assign layer_0[894] = in[157] ^ in[227]; 
    assign layer_0[895] = in[154] ^ in[202]; 
    assign layer_0[896] = in[233] & ~in[166]; 
    assign layer_0[897] = ~(in[115] ^ in[21]); 
    assign layer_0[898] = ~(in[63] ^ in[63]); 
    assign layer_0[899] = ~(in[97] ^ in[98]); 
    assign layer_0[900] = ~(in[181] | in[205]); 
    assign layer_0[901] = in[139] | in[99]; 
    assign layer_0[902] = in[141] ^ in[7]; 
    assign layer_0[903] = in[130] & ~in[188]; 
    assign layer_0[904] = in[126] & ~in[138]; 
    assign layer_0[905] = ~(in[115] | in[243]); 
    assign layer_0[906] = ~in[211] | (in[232] & in[211]); 
    assign layer_0[907] = ~(in[87] ^ in[243]); 
    assign layer_0[908] = ~(in[190] ^ in[65]); 
    assign layer_0[909] = ~in[188] | (in[188] & in[37]); 
    assign layer_0[910] = in[245]; 
    assign layer_0[911] = in[54] & ~in[182]; 
    assign layer_0[912] = in[115] ^ in[113]; 
    assign layer_0[913] = in[183] ^ in[218]; 
    assign layer_0[914] = in[23] ^ in[54]; 
    assign layer_0[915] = ~(in[216] ^ in[247]); 
    assign layer_0[916] = ~(in[152] ^ in[179]); 
    assign layer_0[917] = in[104] & ~in[151]; 
    assign layer_0[918] = ~(in[95] | in[104]); 
    assign layer_0[919] = in[92] ^ in[102]; 
    assign layer_0[920] = in[193] ^ in[157]; 
    assign layer_0[921] = in[9]; 
    assign layer_0[922] = in[152] & ~in[164]; 
    assign layer_0[923] = ~in[214] | (in[214] & in[19]); 
    assign layer_0[924] = in[158]; 
    assign layer_0[925] = in[107] & in[121]; 
    assign layer_0[926] = in[151] ^ in[187]; 
    assign layer_0[927] = ~in[170]; 
    assign layer_0[928] = in[41] & ~in[54]; 
    assign layer_0[929] = ~in[169] | (in[232] & in[169]); 
    assign layer_0[930] = in[85] ^ in[21]; 
    assign layer_0[931] = ~(in[162] ^ in[164]); 
    assign layer_0[932] = in[118] & ~in[162]; 
    assign layer_0[933] = ~(in[179] | in[104]); 
    assign layer_0[934] = ~in[121] | (in[178] & in[121]); 
    assign layer_0[935] = ~(in[227] ^ in[84]); 
    assign layer_0[936] = ~(in[28] | in[194]); 
    assign layer_0[937] = ~(in[34] | in[78]); 
    assign layer_0[938] = in[127] & ~in[219]; 
    assign layer_0[939] = in[56] & ~in[141]; 
    assign layer_0[940] = in[52] ^ in[81]; 
    assign layer_0[941] = in[84] ^ in[71]; 
    assign layer_0[942] = ~(in[116] | in[115]); 
    assign layer_0[943] = ~(in[69] ^ in[38]); 
    assign layer_0[944] = ~in[167]; 
    assign layer_0[945] = in[90] & ~in[196]; 
    assign layer_0[946] = ~in[218] | (in[218] & in[38]); 
    assign layer_0[947] = ~(in[133] ^ in[154]); 
    assign layer_0[948] = in[70]; 
    assign layer_0[949] = ~(in[164] ^ in[183]); 
    assign layer_0[950] = ~(in[185] | in[131]); 
    assign layer_0[951] = in[171] ^ in[125]; 
    assign layer_0[952] = in[55] & ~in[168]; 
    assign layer_0[953] = ~(in[191] ^ in[23]); 
    assign layer_0[954] = ~in[221]; 
    assign layer_0[955] = ~(in[233] ^ in[201]); 
    assign layer_0[956] = ~(in[152] ^ in[8]); 
    assign layer_0[957] = in[77] | in[168]; 
    assign layer_0[958] = in[118] | in[222]; 
    assign layer_0[959] = in[27] | in[7]; 
    assign layer_0[960] = in[7] ^ in[21]; 
    assign layer_0[961] = in[59] & ~in[141]; 
    assign layer_0[962] = in[164] & ~in[246]; 
    assign layer_0[963] = ~(in[182] ^ in[199]); 
    assign layer_0[964] = in[53] & ~in[219]; 
    assign layer_0[965] = in[121]; 
    assign layer_0[966] = in[167] & in[166]; 
    assign layer_0[967] = ~(in[118] ^ in[38]); 
    assign layer_0[968] = ~in[37] | (in[37] & in[171]); 
    assign layer_0[969] = ~in[103]; 
    assign layer_0[970] = in[173] ^ in[196]; 
    assign layer_0[971] = in[92] & ~in[136]; 
    assign layer_0[972] = in[98] & ~in[35]; 
    assign layer_0[973] = in[94] | in[72]; 
    assign layer_0[974] = ~(in[138] ^ in[156]); 
    assign layer_0[975] = ~(in[91] ^ in[71]); 
    assign layer_0[976] = ~(in[190] | in[8]); 
    assign layer_0[977] = in[60] | in[175]; 
    assign layer_0[978] = ~in[135]; 
    assign layer_0[979] = in[212]; 
    assign layer_0[980] = ~(in[219] | in[251]); 
    assign layer_0[981] = in[249] & ~in[167]; 
    assign layer_0[982] = in[142] ^ in[123]; 
    assign layer_0[983] = ~(in[138] ^ in[117]); 
    assign layer_0[984] = in[138] | in[10]; 
    assign layer_0[985] = ~(in[44] | in[123]); 
    assign layer_0[986] = in[60] ^ in[130]; 
    assign layer_0[987] = ~in[89]; 
    assign layer_0[988] = ~(in[87] | in[157]); 
    assign layer_0[989] = in[103] | in[99]; 
    assign layer_0[990] = ~in[9]; 
    assign layer_0[991] = in[8] | in[28]; 
    assign layer_0[992] = ~(in[79] ^ in[124]); 
    assign layer_0[993] = ~(in[133] | in[20]); 
    assign layer_0[994] = in[36] & ~in[67]; 
    assign layer_0[995] = ~(in[164] | in[211]); 
    assign layer_0[996] = in[137] ^ in[55]; 
    assign layer_0[997] = in[231] ^ in[136]; 
    assign layer_0[998] = ~(in[178] ^ in[196]); 
    assign layer_0[999] = in[197] | in[173]; 
    assign layer_0[1000] = ~(in[132] ^ in[10]); 
    assign layer_0[1001] = ~(in[71] ^ in[74]); 
    assign layer_0[1002] = in[59] ^ in[90]; 
    assign layer_0[1003] = in[231] ^ in[250]; 
    assign layer_0[1004] = in[157] | in[35]; 
    assign layer_0[1005] = ~in[168] | (in[69] & in[168]); 
    assign layer_0[1006] = in[99] ^ in[97]; 
    assign layer_0[1007] = ~(in[133] | in[78]); 
    assign layer_0[1008] = in[150] | in[19]; 
    assign layer_0[1009] = ~(in[87] ^ in[57]); 
    assign layer_0[1010] = in[186]; 
    assign layer_0[1011] = ~in[61] | (in[143] & in[61]); 
    assign layer_0[1012] = in[163] ^ in[165]; 
    assign layer_0[1013] = in[47] | in[63]; 
    assign layer_0[1014] = in[8] ^ in[34]; 
    assign layer_0[1015] = ~in[172] | (in[210] & in[172]); 
    assign layer_0[1016] = ~(in[78] | in[83]); 
    assign layer_0[1017] = in[242] | in[80]; 
    assign layer_0[1018] = in[124] | in[110]; 
    assign layer_0[1019] = in[197] | in[161]; 
    assign layer_0[1020] = ~in[47]; 
    assign layer_0[1021] = ~(in[88] ^ in[90]); 
    assign layer_0[1022] = in[40] & ~in[45]; 
    assign layer_0[1023] = ~(in[206] ^ in[197]); 
    assign layer_0[1024] = in[120] & ~in[109]; 
    assign layer_0[1025] = in[58] | in[252]; 
    assign layer_0[1026] = in[75] ^ in[61]; 
    assign layer_0[1027] = ~(in[134] ^ in[40]); 
    assign layer_0[1028] = ~in[101] | (in[101] & in[215]); 
    assign layer_0[1029] = ~(in[101] ^ in[100]); 
    assign layer_0[1030] = in[93] | in[82]; 
    assign layer_0[1031] = in[11] ^ in[29]; 
    assign layer_0[1032] = in[60] ^ in[138]; 
    assign layer_0[1033] = ~(in[99] | in[30]); 
    assign layer_0[1034] = 1'b0; 
    assign layer_0[1035] = ~(in[217] | in[201]); 
    assign layer_0[1036] = in[133] | in[131]; 
    assign layer_0[1037] = in[89] & ~in[184]; 
    assign layer_0[1038] = ~in[92] | (in[92] & in[149]); 
    assign layer_0[1039] = in[179] & in[109]; 
    assign layer_0[1040] = in[172]; 
    assign layer_0[1041] = in[104] | in[135]; 
    assign layer_0[1042] = ~(in[138] ^ in[168]); 
    assign layer_0[1043] = in[95] | in[107]; 
    assign layer_0[1044] = ~in[69]; 
    assign layer_0[1045] = ~in[181] | (in[236] & in[181]); 
    assign layer_0[1046] = in[59] | in[45]; 
    assign layer_0[1047] = in[19] ^ in[155]; 
    assign layer_0[1048] = ~in[46]; 
    assign layer_0[1049] = in[19]; 
    assign layer_0[1050] = ~(in[34] | in[242]); 
    assign layer_0[1051] = in[198] | in[142]; 
    assign layer_0[1052] = in[229] & ~in[198]; 
    assign layer_0[1053] = in[57] & ~in[151]; 
    assign layer_0[1054] = ~(in[79] | in[210]); 
    assign layer_0[1055] = in[63]; 
    assign layer_0[1056] = ~(in[170] ^ in[155]); 
    assign layer_0[1057] = ~(in[171] ^ in[120]); 
    assign layer_0[1058] = ~(in[72] ^ in[38]); 
    assign layer_0[1059] = ~(in[58] | in[42]); 
    assign layer_0[1060] = ~(in[67] | in[69]); 
    assign layer_0[1061] = in[194] ^ in[70]; 
    assign layer_0[1062] = ~in[59] | (in[186] & in[59]); 
    assign layer_0[1063] = ~in[132]; 
    assign layer_0[1064] = ~(in[170] | in[155]); 
    assign layer_0[1065] = ~(in[215] ^ in[171]); 
    assign layer_0[1066] = in[62] | in[158]; 
    assign layer_0[1067] = in[184] | in[162]; 
    assign layer_0[1068] = in[83] ^ in[74]; 
    assign layer_0[1069] = in[42]; 
    assign layer_0[1070] = ~(in[187] ^ in[234]); 
    assign layer_0[1071] = ~(in[241] ^ in[8]); 
    assign layer_0[1072] = ~(in[126] | in[214]); 
    assign layer_0[1073] = ~in[104] | (in[104] & in[148]); 
    assign layer_0[1074] = in[146] ^ in[121]; 
    assign layer_0[1075] = in[8] | in[6]; 
    assign layer_0[1076] = ~in[76] | (in[76] & in[29]); 
    assign layer_0[1077] = ~in[139]; 
    assign layer_0[1078] = ~in[197] | (in[197] & in[188]); 
    assign layer_0[1079] = ~(in[52] | in[42]); 
    assign layer_0[1080] = in[229] | in[53]; 
    assign layer_0[1081] = in[100] ^ in[47]; 
    assign layer_0[1082] = ~in[165]; 
    assign layer_0[1083] = ~(in[245] ^ in[217]); 
    assign layer_0[1084] = in[119]; 
    assign layer_0[1085] = in[46] ^ in[79]; 
    assign layer_0[1086] = ~(in[24] | in[158]); 
    assign layer_0[1087] = in[214] ^ in[58]; 
    assign layer_0[1088] = ~(in[183] ^ in[135]); 
    assign layer_0[1089] = ~in[182] | (in[182] & in[90]); 
    assign layer_0[1090] = in[68] ^ in[42]; 
    assign layer_0[1091] = ~in[35] | (in[35] & in[30]); 
    assign layer_0[1092] = in[9] | in[21]; 
    assign layer_0[1093] = in[124] ^ in[83]; 
    assign layer_0[1094] = ~(in[132] ^ in[147]); 
    assign layer_0[1095] = in[167]; 
    assign layer_0[1096] = in[139] ^ in[171]; 
    assign layer_0[1097] = in[52]; 
    assign layer_0[1098] = in[229]; 
    assign layer_0[1099] = ~(in[203] ^ in[248]); 
    assign layer_0[1100] = in[20] | in[210]; 
    assign layer_0[1101] = ~in[90] | (in[232] & in[90]); 
    assign layer_0[1102] = in[124]; 
    assign layer_0[1103] = ~(in[75] ^ in[77]); 
    assign layer_0[1104] = in[185] ^ in[218]; 
    assign layer_0[1105] = in[135] ^ in[151]; 
    assign layer_0[1106] = in[100] ^ in[87]; 
    assign layer_0[1107] = in[153] & ~in[102]; 
    assign layer_0[1108] = ~in[217] | (in[214] & in[217]); 
    assign layer_0[1109] = ~(in[219] ^ in[58]); 
    assign layer_0[1110] = ~(in[229] | in[228]); 
    assign layer_0[1111] = ~in[38]; 
    assign layer_0[1112] = in[86] ^ in[41]; 
    assign layer_0[1113] = in[66] ^ in[150]; 
    assign layer_0[1114] = in[122] & in[106]; 
    assign layer_0[1115] = ~(in[219] | in[187]); 
    assign layer_0[1116] = in[101] & ~in[22]; 
    assign layer_0[1117] = ~(in[178] ^ in[65]); 
    assign layer_0[1118] = in[46] ^ in[94]; 
    assign layer_0[1119] = ~(in[84] | in[221]); 
    assign layer_0[1120] = ~(in[149] | in[229]); 
    assign layer_0[1121] = in[231] ^ in[183]; 
    assign layer_0[1122] = in[214] ^ in[245]; 
    assign layer_0[1123] = ~(in[244] ^ in[124]); 
    assign layer_0[1124] = ~(in[102] ^ in[87]); 
    assign layer_0[1125] = ~(in[165] ^ in[148]); 
    assign layer_0[1126] = in[57] | in[81]; 
    assign layer_0[1127] = in[100] ^ in[102]; 
    assign layer_0[1128] = ~(in[137] ^ in[172]); 
    assign layer_0[1129] = in[38] ^ in[234]; 
    assign layer_0[1130] = in[45] ^ in[79]; 
    assign layer_0[1131] = ~in[194]; 
    assign layer_0[1132] = ~(in[198] ^ in[244]); 
    assign layer_0[1133] = ~in[130]; 
    assign layer_0[1134] = ~(in[203] | in[29]); 
    assign layer_0[1135] = ~(in[204] ^ in[193]); 
    assign layer_0[1136] = in[148] | in[246]; 
    assign layer_0[1137] = ~(in[190] ^ in[7]); 
    assign layer_0[1138] = ~(in[214] ^ in[22]); 
    assign layer_0[1139] = ~(in[77] | in[78]); 
    assign layer_0[1140] = 1'b0; 
    assign layer_0[1141] = ~(in[59] & in[77]); 
    assign layer_0[1142] = in[151] ^ in[198]; 
    assign layer_0[1143] = ~(in[37] ^ in[186]); 
    assign layer_0[1144] = ~(in[236] | in[86]); 
    assign layer_0[1145] = ~(in[186] ^ in[234]); 
    assign layer_0[1146] = ~(in[78] | in[53]); 
    assign layer_0[1147] = ~(in[52] | in[207]); 
    assign layer_0[1148] = ~(in[160] ^ in[34]); 
    assign layer_0[1149] = ~(in[152] | in[140]); 
    assign layer_0[1150] = ~(in[182] | in[104]); 
    assign layer_0[1151] = in[235] ^ in[221]; 
    assign layer_0[1152] = ~(in[50] | in[186]); 
    assign layer_0[1153] = ~(in[231] ^ in[134]); 
    assign layer_0[1154] = ~(in[132] ^ in[150]); 
    assign layer_0[1155] = ~(in[218] ^ in[220]); 
    assign layer_0[1156] = ~in[9] | (in[171] & in[9]); 
    assign layer_0[1157] = ~(in[197] | in[127]); 
    assign layer_0[1158] = ~in[133]; 
    assign layer_0[1159] = ~(in[216] | in[189]); 
    assign layer_0[1160] = in[107] ^ in[156]; 
    assign layer_0[1161] = in[72]; 
    assign layer_0[1162] = in[71] ^ in[39]; 
    assign layer_0[1163] = in[20]; 
    assign layer_0[1164] = in[248] | in[200]; 
    assign layer_0[1165] = in[135]; 
    assign layer_0[1166] = ~in[179] | (in[179] & in[121]); 
    assign layer_0[1167] = ~(in[148] ^ in[212]); 
    assign layer_0[1168] = ~in[198] | (in[198] & in[12]); 
    assign layer_0[1169] = ~(in[215] ^ in[162]); 
    assign layer_0[1170] = in[182] ^ in[164]; 
    assign layer_0[1171] = 1'b1; 
    assign layer_0[1172] = in[134] & ~in[59]; 
    assign layer_0[1173] = ~(in[241] | in[100]); 
    assign layer_0[1174] = ~(in[94] ^ in[184]); 
    assign layer_0[1175] = ~(in[201] ^ in[105]); 
    assign layer_0[1176] = ~(in[164] | in[183]); 
    assign layer_0[1177] = ~in[182]; 
    assign layer_0[1178] = in[38]; 
    assign layer_0[1179] = in[73] ^ in[88]; 
    assign layer_0[1180] = ~(in[119] ^ in[148]); 
    assign layer_0[1181] = in[51] ^ in[155]; 
    assign layer_0[1182] = ~(in[155] | in[243]); 
    assign layer_0[1183] = in[184] ^ in[67]; 
    assign layer_0[1184] = ~(in[213] ^ in[61]); 
    assign layer_0[1185] = in[218] | in[140]; 
    assign layer_0[1186] = in[44] | in[39]; 
    assign layer_0[1187] = ~(in[107] ^ in[139]); 
    assign layer_0[1188] = ~(in[119] ^ in[149]); 
    assign layer_0[1189] = ~(in[51] | in[213]); 
    assign layer_0[1190] = in[242] ^ in[99]; 
    assign layer_0[1191] = ~(in[120] ^ in[104]); 
    assign layer_0[1192] = ~(in[139] ^ in[141]); 
    assign layer_0[1193] = in[239] | in[252]; 
    assign layer_0[1194] = in[76] | in[40]; 
    assign layer_0[1195] = ~(in[249] | in[236]); 
    assign layer_0[1196] = in[213] ^ in[78]; 
    assign layer_0[1197] = ~in[188] | (in[188] & in[129]); 
    assign layer_0[1198] = in[91] ^ in[93]; 
    assign layer_0[1199] = in[100] ^ in[182]; 
    assign layer_0[1200] = in[10] ^ in[20]; 
    assign layer_0[1201] = in[38]; 
    assign layer_0[1202] = ~in[179] | (in[179] & in[47]); 
    assign layer_0[1203] = ~(in[148] | in[123]); 
    assign layer_0[1204] = in[231] & ~in[152]; 
    assign layer_0[1205] = ~(in[114] | in[226]); 
    assign layer_0[1206] = in[90] & ~in[196]; 
    assign layer_0[1207] = ~in[87]; 
    assign layer_0[1208] = in[57] ^ in[141]; 
    assign layer_0[1209] = ~in[36] | (in[36] & in[215]); 
    assign layer_0[1210] = ~(in[73] ^ in[38]); 
    assign layer_0[1211] = in[57] ^ in[88]; 
    assign layer_0[1212] = ~in[51] | (in[227] & in[51]); 
    assign layer_0[1213] = in[23] | in[187]; 
    assign layer_0[1214] = ~(in[40] ^ in[98]); 
    assign layer_0[1215] = ~in[155] | (in[210] & in[155]); 
    assign layer_0[1216] = ~in[56]; 
    assign layer_0[1217] = ~(in[73] & in[214]); 
    assign layer_0[1218] = ~(in[123] ^ in[76]); 
    assign layer_0[1219] = in[133] & ~in[136]; 
    assign layer_0[1220] = in[118] | in[210]; 
    assign layer_0[1221] = ~(in[180] | in[194]); 
    assign layer_0[1222] = in[67] ^ in[104]; 
    assign layer_0[1223] = ~(in[149] ^ in[127]); 
    assign layer_0[1224] = ~(in[66] ^ in[35]); 
    assign layer_0[1225] = in[111] ^ in[109]; 
    assign layer_0[1226] = ~in[209] | (in[117] & in[209]); 
    assign layer_0[1227] = ~in[115] | (in[115] & in[192]); 
    assign layer_0[1228] = ~(in[99] | in[87]); 
    assign layer_0[1229] = ~in[88]; 
    assign layer_0[1230] = ~(in[135] | in[195]); 
    assign layer_0[1231] = in[166] ^ in[211]; 
    assign layer_0[1232] = ~(in[11] | in[102]); 
    assign layer_0[1233] = in[220] ^ in[250]; 
    assign layer_0[1234] = in[244] ^ in[83]; 
    assign layer_0[1235] = in[77] ^ in[139]; 
    assign layer_0[1236] = in[107] ^ in[118]; 
    assign layer_0[1237] = ~in[24] | (in[24] & in[42]); 
    assign layer_0[1238] = in[164]; 
    assign layer_0[1239] = in[168]; 
    assign layer_0[1240] = ~(in[60] ^ in[234]); 
    assign layer_0[1241] = ~(in[55] & in[69]); 
    assign layer_0[1242] = ~(in[196] ^ in[204]); 
    assign layer_0[1243] = ~(in[152] ^ in[121]); 
    assign layer_0[1244] = in[83] | in[120]; 
    assign layer_0[1245] = in[149] ^ in[147]; 
    assign layer_0[1246] = ~(in[179] ^ in[236]); 
    assign layer_0[1247] = ~(in[181] ^ in[78]); 
    assign layer_0[1248] = ~(in[88] ^ in[120]); 
    assign layer_0[1249] = in[197]; 
    assign layer_0[1250] = in[182] & ~in[116]; 
    assign layer_0[1251] = in[186] | in[85]; 
    assign layer_0[1252] = in[90] | in[105]; 
    assign layer_0[1253] = ~in[122] | (in[122] & in[172]); 
    assign layer_0[1254] = ~(in[220] | in[23]); 
    assign layer_0[1255] = in[111] ^ in[109]; 
    assign layer_0[1256] = ~(in[188] ^ in[154]); 
    assign layer_0[1257] = ~(in[78] | in[77]); 
    assign layer_0[1258] = in[124] ^ in[252]; 
    assign layer_0[1259] = in[221] ^ in[111]; 
    assign layer_0[1260] = ~(in[53] ^ in[134]); 
    assign layer_0[1261] = ~in[120] | (in[138] & in[120]); 
    assign layer_0[1262] = 1'b1; 
    assign layer_0[1263] = in[60] ^ in[166]; 
    assign layer_0[1264] = ~in[36]; 
    assign layer_0[1265] = ~in[199] | (in[109] & in[199]); 
    assign layer_0[1266] = ~(in[84] ^ in[119]); 
    assign layer_0[1267] = in[176]; 
    assign layer_0[1268] = ~(in[124] | in[58]); 
    assign layer_0[1269] = ~(in[135] ^ in[103]); 
    assign layer_0[1270] = in[30]; 
    assign layer_0[1271] = ~in[231] | (in[231] & in[76]); 
    assign layer_0[1272] = in[59] | in[61]; 
    assign layer_0[1273] = in[148] | in[220]; 
    assign layer_0[1274] = ~(in[157] ^ in[193]); 
    assign layer_0[1275] = ~(in[190] ^ in[225]); 
    assign layer_0[1276] = ~(in[147] ^ in[120]); 
    assign layer_0[1277] = in[110] | in[155]; 
    assign layer_0[1278] = ~in[70] | (in[164] & in[70]); 
    assign layer_0[1279] = in[231] & ~in[107]; 
    assign layer_0[1280] = in[68] ^ in[85]; 
    assign layer_0[1281] = in[21] ^ in[91]; 
    assign layer_0[1282] = ~in[218] | (in[218] & in[81]); 
    assign layer_0[1283] = ~(in[101] ^ in[170]); 
    assign layer_0[1284] = ~(in[98] ^ in[169]); 
    assign layer_0[1285] = ~(in[62] ^ in[73]); 
    assign layer_0[1286] = in[138] | in[197]; 
    assign layer_0[1287] = ~in[121] | (in[181] & in[121]); 
    assign layer_0[1288] = in[107] & in[120]; 
    assign layer_0[1289] = in[230]; 
    assign layer_0[1290] = in[86] ^ in[120]; 
    assign layer_0[1291] = in[118] & ~in[105]; 
    assign layer_0[1292] = ~in[136] | (in[187] & in[136]); 
    assign layer_0[1293] = in[244] ^ in[195]; 
    assign layer_0[1294] = in[62] | in[68]; 
    assign layer_0[1295] = ~in[26] | (in[26] & in[245]); 
    assign layer_0[1296] = ~(in[79] ^ in[51]); 
    assign layer_0[1297] = in[19] ^ in[76]; 
    assign layer_0[1298] = ~(in[39] ^ in[122]); 
    assign layer_0[1299] = ~(in[102] | in[101]); 
    assign layer_0[1300] = ~(in[88] ^ in[214]); 
    assign layer_0[1301] = in[119] ^ in[113]; 
    assign layer_0[1302] = in[115] | in[200]; 
    assign layer_0[1303] = in[214] ^ in[199]; 
    assign layer_0[1304] = ~in[183] | (in[183] & in[249]); 
    assign layer_0[1305] = ~in[132] | (in[11] & in[132]); 
    assign layer_0[1306] = in[105] ^ in[107]; 
    assign layer_0[1307] = ~(in[93] ^ in[110]); 
    assign layer_0[1308] = in[88] ^ in[119]; 
    assign layer_0[1309] = in[102] ^ in[70]; 
    assign layer_0[1310] = in[7] ^ in[143]; 
    assign layer_0[1311] = in[141]; 
    assign layer_0[1312] = ~in[104] | (in[123] & in[104]); 
    assign layer_0[1313] = in[92] ^ in[199]; 
    assign layer_0[1314] = ~(in[177] | in[155]); 
    assign layer_0[1315] = ~in[105]; 
    assign layer_0[1316] = in[169] | in[57]; 
    assign layer_0[1317] = in[138]; 
    assign layer_0[1318] = in[38] & ~in[19]; 
    assign layer_0[1319] = ~(in[218] ^ in[186]); 
    assign layer_0[1320] = ~(in[159] ^ in[28]); 
    assign layer_0[1321] = in[210] | in[251]; 
    assign layer_0[1322] = ~(in[170] | in[142]); 
    assign layer_0[1323] = in[5] | in[127]; 
    assign layer_0[1324] = in[212] ^ in[71]; 
    assign layer_0[1325] = ~in[166] | (in[214] & in[166]); 
    assign layer_0[1326] = ~(in[30] ^ in[93]); 
    assign layer_0[1327] = in[182] & ~in[78]; 
    assign layer_0[1328] = ~(in[153] ^ in[156]); 
    assign layer_0[1329] = ~(in[140] ^ in[183]); 
    assign layer_0[1330] = ~(in[198] ^ in[180]); 
    assign layer_0[1331] = ~(in[76] ^ in[78]); 
    assign layer_0[1332] = ~(in[229] | in[227]); 
    assign layer_0[1333] = in[44] | in[61]; 
    assign layer_0[1334] = in[246]; 
    assign layer_0[1335] = ~(in[150] ^ in[25]); 
    assign layer_0[1336] = ~(in[76] | in[90]); 
    assign layer_0[1337] = in[232] ^ in[153]; 
    assign layer_0[1338] = in[119] | in[77]; 
    assign layer_0[1339] = in[105] & ~in[152]; 
    assign layer_0[1340] = ~(in[54] | in[99]); 
    assign layer_0[1341] = in[239] | in[107]; 
    assign layer_0[1342] = in[9] & ~in[102]; 
    assign layer_0[1343] = ~in[191]; 
    assign layer_0[1344] = ~(in[166] | in[174]); 
    assign layer_0[1345] = in[73] | in[58]; 
    assign layer_0[1346] = ~(in[167] ^ in[165]); 
    assign layer_0[1347] = in[179] ^ in[197]; 
    assign layer_0[1348] = in[244] | in[165]; 
    assign layer_0[1349] = ~(in[218] ^ in[212]); 
    assign layer_0[1350] = ~(in[166] ^ in[164]); 
    assign layer_0[1351] = ~in[56] | (in[203] & in[56]); 
    assign layer_0[1352] = ~in[116] | (in[186] & in[116]); 
    assign layer_0[1353] = in[53] ^ in[101]; 
    assign layer_0[1354] = in[116] ^ in[150]; 
    assign layer_0[1355] = ~(in[134] | in[170]); 
    assign layer_0[1356] = ~(in[119] ^ in[150]); 
    assign layer_0[1357] = ~in[179]; 
    assign layer_0[1358] = in[25] ^ in[58]; 
    assign layer_0[1359] = ~(in[104] | in[133]); 
    assign layer_0[1360] = in[182] ^ in[220]; 
    assign layer_0[1361] = in[40] ^ in[87]; 
    assign layer_0[1362] = ~(in[59] | in[124]); 
    assign layer_0[1363] = ~in[104] | (in[139] & in[104]); 
    assign layer_0[1364] = in[165] ^ in[8]; 
    assign layer_0[1365] = ~(in[216] ^ in[234]); 
    assign layer_0[1366] = ~in[252]; 
    assign layer_0[1367] = in[85] ^ in[87]; 
    assign layer_0[1368] = in[81]; 
    assign layer_0[1369] = in[163] | in[182]; 
    assign layer_0[1370] = in[100]; 
    assign layer_0[1371] = in[85] ^ in[52]; 
    assign layer_0[1372] = in[89] & ~in[104]; 
    assign layer_0[1373] = ~(in[220] | in[222]); 
    assign layer_0[1374] = ~(in[85] | in[252]); 
    assign layer_0[1375] = ~(in[159] | in[89]); 
    assign layer_0[1376] = ~(in[187] | in[157]); 
    assign layer_0[1377] = ~(in[178] ^ in[107]); 
    assign layer_0[1378] = in[185]; 
    assign layer_0[1379] = in[36] ^ in[235]; 
    assign layer_0[1380] = 1'b1; 
    assign layer_0[1381] = ~(in[134] | in[150]); 
    assign layer_0[1382] = ~in[74] | (in[74] & in[46]); 
    assign layer_0[1383] = ~in[50] | (in[110] & in[50]); 
    assign layer_0[1384] = ~in[42] | (in[248] & in[42]); 
    assign layer_0[1385] = in[74] & ~in[61]; 
    assign layer_0[1386] = in[185] ^ in[211]; 
    assign layer_0[1387] = ~(in[70] ^ in[23]); 
    assign layer_0[1388] = ~in[74] | (in[74] & in[251]); 
    assign layer_0[1389] = ~in[149] | (in[53] & in[149]); 
    assign layer_0[1390] = ~(in[183] ^ in[165]); 
    assign layer_0[1391] = in[179] & in[30]; 
    assign layer_0[1392] = in[103] ^ in[117]; 
    assign layer_0[1393] = ~in[245]; 
    assign layer_0[1394] = in[99] | in[248]; 
    assign layer_0[1395] = in[181] ^ in[230]; 
    assign layer_0[1396] = ~(in[58] ^ in[89]); 
    assign layer_0[1397] = ~(in[177] | in[67]); 
    assign layer_0[1398] = ~in[182] | (in[57] & in[182]); 
    assign layer_0[1399] = ~(in[78] ^ in[104]); 
    assign layer_0[1400] = in[89] ^ in[107]; 
    assign layer_0[1401] = ~(in[149] | in[244]); 
    assign layer_0[1402] = ~(in[110] | in[85]); 
    assign layer_0[1403] = ~(in[206] ^ in[174]); 
    assign layer_0[1404] = ~in[41] | (in[123] & in[41]); 
    assign layer_0[1405] = in[132] & in[148]; 
    assign layer_0[1406] = ~(in[36] | in[101]); 
    assign layer_0[1407] = ~(in[107] ^ in[94]); 
    assign layer_0[1408] = in[79] ^ in[228]; 
    assign layer_0[1409] = ~(in[57] | in[104]); 
    assign layer_0[1410] = ~(in[165] ^ in[147]); 
    assign layer_0[1411] = ~(in[134] | in[21]); 
    assign layer_0[1412] = in[119] ^ in[102]; 
    assign layer_0[1413] = in[135] | in[194]; 
    assign layer_0[1414] = in[227] ^ in[136]; 
    assign layer_0[1415] = ~(in[81] | in[50]); 
    assign layer_0[1416] = ~(in[196] ^ in[182]); 
    assign layer_0[1417] = ~(in[42] ^ in[76]); 
    assign layer_0[1418] = ~(in[132] | in[130]); 
    assign layer_0[1419] = in[132] & ~in[183]; 
    assign layer_0[1420] = ~(in[137] ^ in[171]); 
    assign layer_0[1421] = 1'b0; 
    assign layer_0[1422] = in[72] ^ in[44]; 
    assign layer_0[1423] = in[167] | in[79]; 
    assign layer_0[1424] = ~in[42]; 
    assign layer_0[1425] = ~in[115]; 
    assign layer_0[1426] = in[154] & ~in[194]; 
    assign layer_0[1427] = ~(in[79] ^ in[114]); 
    assign layer_0[1428] = in[46] ^ in[63]; 
    assign layer_0[1429] = ~(in[163] | in[75]); 
    assign layer_0[1430] = ~(in[193] | in[135]); 
    assign layer_0[1431] = ~(in[23] ^ in[163]); 
    assign layer_0[1432] = in[42] ^ in[89]; 
    assign layer_0[1433] = in[108] ^ in[94]; 
    assign layer_0[1434] = in[183]; 
    assign layer_0[1435] = in[36] | in[179]; 
    assign layer_0[1436] = ~in[218]; 
    assign layer_0[1437] = in[173] ^ in[111]; 
    assign layer_0[1438] = ~in[154]; 
    assign layer_0[1439] = in[36] & ~in[68]; 
    assign layer_0[1440] = in[106] ^ in[95]; 
    assign layer_0[1441] = ~(in[108] ^ in[232]); 
    assign layer_0[1442] = in[124] ^ in[92]; 
    assign layer_0[1443] = in[107] ^ in[23]; 
    assign layer_0[1444] = in[63] | in[54]; 
    assign layer_0[1445] = ~(in[166] ^ in[230]); 
    assign layer_0[1446] = in[166] | in[149]; 
    assign layer_0[1447] = in[124]; 
    assign layer_0[1448] = in[85] ^ in[24]; 
    assign layer_0[1449] = in[105] ^ in[10]; 
    assign layer_0[1450] = in[231] | in[244]; 
    assign layer_0[1451] = ~(in[135] & in[136]); 
    assign layer_0[1452] = in[220]; 
    assign layer_0[1453] = in[155]; 
    assign layer_0[1454] = in[235] | in[152]; 
    assign layer_0[1455] = ~(in[131] ^ in[129]); 
    assign layer_0[1456] = ~in[188]; 
    assign layer_0[1457] = in[137] ^ in[146]; 
    assign layer_0[1458] = ~in[152] | (in[152] & in[146]); 
    assign layer_0[1459] = in[71] & ~in[179]; 
    assign layer_0[1460] = ~(in[179] | in[200]); 
    assign layer_0[1461] = in[22] | in[37]; 
    assign layer_0[1462] = ~(in[84] ^ in[98]); 
    assign layer_0[1463] = in[93] ^ in[171]; 
    assign layer_0[1464] = in[115] ^ in[113]; 
    assign layer_0[1465] = in[103]; 
    assign layer_0[1466] = in[72] | in[112]; 
    assign layer_0[1467] = in[109] ^ in[106]; 
    assign layer_0[1468] = ~(in[211] | in[165]); 
    assign layer_0[1469] = ~(in[135] ^ in[152]); 
    assign layer_0[1470] = ~(in[140] ^ in[122]); 
    assign layer_0[1471] = in[142] & ~in[138]; 
    assign layer_0[1472] = ~(in[73] ^ in[97]); 
    assign layer_0[1473] = in[169] & ~in[214]; 
    assign layer_0[1474] = ~(in[37] | in[27]); 
    assign layer_0[1475] = ~(in[176] | in[176]); 
    assign layer_0[1476] = ~(in[153] ^ in[119]); 
    assign layer_0[1477] = ~(in[152] | in[137]); 
    assign layer_0[1478] = ~(in[39] ^ in[76]); 
    assign layer_0[1479] = ~(in[134] ^ in[164]); 
    assign layer_0[1480] = ~(in[85] ^ in[100]); 
    assign layer_0[1481] = ~(in[166] | in[211]); 
    assign layer_0[1482] = in[232] & ~in[106]; 
    assign layer_0[1483] = in[93] | in[151]; 
    assign layer_0[1484] = ~(in[202] & in[156]); 
    assign layer_0[1485] = in[196] ^ in[237]; 
    assign layer_0[1486] = ~in[147]; 
    assign layer_0[1487] = in[63] | in[30]; 
    assign layer_0[1488] = in[91] ^ in[89]; 
    assign layer_0[1489] = ~(in[99] ^ in[102]); 
    assign layer_0[1490] = ~in[218] | (in[101] & in[218]); 
    assign layer_0[1491] = ~(in[108] ^ in[61]); 
    assign layer_0[1492] = ~(in[56] ^ in[25]); 
    assign layer_0[1493] = in[159] ^ in[12]; 
    assign layer_0[1494] = ~(in[197] ^ in[231]); 
    assign layer_0[1495] = in[211] ^ in[72]; 
    assign layer_0[1496] = ~(in[149] ^ in[163]); 
    assign layer_0[1497] = ~(in[88] ^ in[44]); 
    assign layer_0[1498] = ~in[184]; 
    assign layer_0[1499] = ~(in[204] ^ in[235]); 
    assign layer_0[1500] = ~in[162]; 
    assign layer_0[1501] = ~in[19]; 
    assign layer_0[1502] = in[78]; 
    assign layer_0[1503] = ~(in[93] ^ in[91]); 
    assign layer_0[1504] = in[28] | in[143]; 
    assign layer_0[1505] = ~in[10] | (in[37] & in[10]); 
    assign layer_0[1506] = ~in[115]; 
    assign layer_0[1507] = in[108] ^ in[91]; 
    assign layer_0[1508] = in[190] ^ in[95]; 
    assign layer_0[1509] = in[70] ^ in[38]; 
    assign layer_0[1510] = in[131] & ~in[179]; 
    assign layer_0[1511] = ~in[197]; 
    assign layer_0[1512] = ~(in[103] | in[99]); 
    assign layer_0[1513] = ~in[36]; 
    assign layer_0[1514] = ~(in[77] | in[247]); 
    assign layer_0[1515] = ~(in[117] | in[131]); 
    assign layer_0[1516] = in[174]; 
    assign layer_0[1517] = ~in[108] | (in[95] & in[108]); 
    assign layer_0[1518] = in[166] ^ in[135]; 
    assign layer_0[1519] = ~(in[100] ^ in[86]); 
    assign layer_0[1520] = in[93] ^ in[45]; 
    assign layer_0[1521] = in[155] | in[123]; 
    assign layer_0[1522] = in[121] & ~in[139]; 
    assign layer_0[1523] = ~in[88] | (in[88] & in[42]); 
    assign layer_0[1524] = in[196] ^ in[62]; 
    assign layer_0[1525] = ~in[247]; 
    assign layer_0[1526] = in[34] ^ in[162]; 
    assign layer_0[1527] = in[220] | in[205]; 
    assign layer_0[1528] = ~(in[108] ^ in[167]); 
    assign layer_0[1529] = ~(in[34] | in[147]); 
    assign layer_0[1530] = ~in[100] | (in[100] & in[24]); 
    assign layer_0[1531] = in[187] ^ in[218]; 
    assign layer_0[1532] = in[107] | in[150]; 
    assign layer_0[1533] = in[102] ^ in[53]; 
    assign layer_0[1534] = in[166] ^ in[135]; 
    assign layer_0[1535] = in[136] ^ in[105]; 
    assign layer_0[1536] = in[137] & ~in[156]; 
    assign layer_0[1537] = in[81] | in[52]; 
    assign layer_0[1538] = in[22] | in[20]; 
    assign layer_0[1539] = ~(in[126] ^ in[74]); 
    assign layer_0[1540] = in[190] | in[158]; 
    assign layer_0[1541] = ~(in[230] ^ in[98]); 
    assign layer_0[1542] = ~(in[8] ^ in[147]); 
    assign layer_0[1543] = ~(in[49] | in[94]); 
    assign layer_0[1544] = in[56] & ~in[147]; 
    assign layer_0[1545] = ~(in[87] ^ in[42]); 
    assign layer_0[1546] = ~(in[178] | in[180]); 
    assign layer_0[1547] = in[201] | in[232]; 
    assign layer_0[1548] = ~(in[121] ^ in[167]); 
    assign layer_0[1549] = in[236] ^ in[220]; 
    assign layer_0[1550] = ~(in[101] ^ in[19]); 
    assign layer_0[1551] = in[203]; 
    assign layer_0[1552] = ~(in[162] ^ in[180]); 
    assign layer_0[1553] = in[148] & ~in[66]; 
    assign layer_0[1554] = ~(in[121] ^ in[116]); 
    assign layer_0[1555] = ~(in[29] & in[196]); 
    assign layer_0[1556] = in[89] ^ in[77]; 
    assign layer_0[1557] = ~(in[229] ^ in[196]); 
    assign layer_0[1558] = in[211]; 
    assign layer_0[1559] = in[249] | in[92]; 
    assign layer_0[1560] = ~(in[30] | in[166]); 
    assign layer_0[1561] = ~in[130] | (in[130] & in[120]); 
    assign layer_0[1562] = ~(in[206] ^ in[235]); 
    assign layer_0[1563] = in[229] | in[72]; 
    assign layer_0[1564] = in[73] & ~in[9]; 
    assign layer_0[1565] = ~in[186] | (in[186] & in[210]); 
    assign layer_0[1566] = in[98]; 
    assign layer_0[1567] = ~(in[188] ^ in[219]); 
    assign layer_0[1568] = ~(in[21] | in[237]); 
    assign layer_0[1569] = in[9] | in[27]; 
    assign layer_0[1570] = ~(in[169] ^ in[187]); 
    assign layer_0[1571] = in[219] | in[172]; 
    assign layer_0[1572] = ~(in[177] | in[226]); 
    assign layer_0[1573] = in[72] & ~in[151]; 
    assign layer_0[1574] = ~in[83]; 
    assign layer_0[1575] = ~in[107] | (in[73] & in[107]); 
    assign layer_0[1576] = ~(in[202] ^ in[233]); 
    assign layer_0[1577] = in[90] & ~in[78]; 
    assign layer_0[1578] = in[21] | in[77]; 
    assign layer_0[1579] = in[59] ^ in[89]; 
    assign layer_0[1580] = in[230] | in[151]; 
    assign layer_0[1581] = ~(in[188] ^ in[220]); 
    assign layer_0[1582] = ~(in[36] | in[79]); 
    assign layer_0[1583] = in[21] | in[190]; 
    assign layer_0[1584] = in[158] | in[197]; 
    assign layer_0[1585] = in[104]; 
    assign layer_0[1586] = ~(in[101] ^ in[136]); 
    assign layer_0[1587] = in[120] ^ in[151]; 
    assign layer_0[1588] = ~(in[181] ^ in[202]); 
    assign layer_0[1589] = ~(in[90] ^ in[54]); 
    assign layer_0[1590] = ~(in[60] ^ in[164]); 
    assign layer_0[1591] = ~(in[41] ^ in[43]); 
    assign layer_0[1592] = ~(in[30] | in[149]); 
    assign layer_0[1593] = ~in[136] | (in[136] & in[177]); 
    assign layer_0[1594] = in[181] | in[195]; 
    assign layer_0[1595] = ~(in[9] ^ in[168]); 
    assign layer_0[1596] = ~(in[142] ^ in[88]); 
    assign layer_0[1597] = ~(in[116] ^ in[114]); 
    assign layer_0[1598] = ~(in[55] ^ in[87]); 
    assign layer_0[1599] = ~in[153] | (in[153] & in[235]); 
    assign layer_0[1600] = ~(in[234] | in[213]); 
    assign layer_0[1601] = ~(in[25] | in[38]); 
    assign layer_0[1602] = in[75] | in[249]; 
    assign layer_0[1603] = in[177]; 
    assign layer_0[1604] = ~(in[207] | in[11]); 
    assign layer_0[1605] = in[136] | in[120]; 
    assign layer_0[1606] = ~(in[92] ^ in[55]); 
    assign layer_0[1607] = ~(in[58] ^ in[181]); 
    assign layer_0[1608] = ~(in[133] ^ in[162]); 
    assign layer_0[1609] = ~(in[159] | in[206]); 
    assign layer_0[1610] = ~(in[127] ^ in[9]); 
    assign layer_0[1611] = ~(in[136] ^ in[101]); 
    assign layer_0[1612] = ~(in[99] ^ in[37]); 
    assign layer_0[1613] = ~in[55] | (in[55] & in[186]); 
    assign layer_0[1614] = ~(in[130] ^ in[172]); 
    assign layer_0[1615] = ~in[245]; 
    assign layer_0[1616] = in[181] | in[230]; 
    assign layer_0[1617] = in[107] ^ in[121]; 
    assign layer_0[1618] = in[153] ^ in[133]; 
    assign layer_0[1619] = ~in[102] | (in[84] & in[102]); 
    assign layer_0[1620] = in[163] | in[99]; 
    assign layer_0[1621] = in[167] & ~in[248]; 
    assign layer_0[1622] = in[65]; 
    assign layer_0[1623] = in[10] ^ in[7]; 
    assign layer_0[1624] = ~(in[174] | in[126]); 
    assign layer_0[1625] = in[168] & ~in[212]; 
    assign layer_0[1626] = ~(in[104] | in[97]); 
    assign layer_0[1627] = in[228] | in[243]; 
    assign layer_0[1628] = ~(in[102] ^ in[54]); 
    assign layer_0[1629] = ~(in[155] | in[195]); 
    assign layer_0[1630] = ~(in[77] | in[62]); 
    assign layer_0[1631] = in[41] & ~in[109]; 
    assign layer_0[1632] = in[54] ^ in[109]; 
    assign layer_0[1633] = in[73] | in[95]; 
    assign layer_0[1634] = ~(in[232] ^ in[25]); 
    assign layer_0[1635] = in[124]; 
    assign layer_0[1636] = ~(in[245] ^ in[229]); 
    assign layer_0[1637] = in[58] & ~in[181]; 
    assign layer_0[1638] = ~(in[184] ^ in[149]); 
    assign layer_0[1639] = in[88] & ~in[107]; 
    assign layer_0[1640] = in[250] ^ in[122]; 
    assign layer_0[1641] = ~(in[76] ^ in[74]); 
    assign layer_0[1642] = in[134] & ~in[116]; 
    assign layer_0[1643] = in[106] ^ in[108]; 
    assign layer_0[1644] = in[5] ^ in[179]; 
    assign layer_0[1645] = ~(in[196] ^ in[203]); 
    assign layer_0[1646] = ~in[100] | (in[100] & in[132]); 
    assign layer_0[1647] = in[213] ^ in[134]; 
    assign layer_0[1648] = in[103] & ~in[54]; 
    assign layer_0[1649] = ~(in[84] ^ in[98]); 
    assign layer_0[1650] = in[247] ^ in[243]; 
    assign layer_0[1651] = in[228] & ~in[140]; 
    assign layer_0[1652] = ~in[150] | (in[150] & in[105]); 
    assign layer_0[1653] = in[136] ^ in[167]; 
    assign layer_0[1654] = in[143]; 
    assign layer_0[1655] = in[168]; 
    assign layer_0[1656] = in[118] ^ in[116]; 
    assign layer_0[1657] = in[186] ^ in[34]; 
    assign layer_0[1658] = ~in[98]; 
    assign layer_0[1659] = ~in[92]; 
    assign layer_0[1660] = in[209] ^ in[11]; 
    assign layer_0[1661] = ~in[199] | (in[199] & in[148]); 
    assign layer_0[1662] = ~(in[52] & in[185]); 
    assign layer_0[1663] = in[251] | in[244]; 
    assign layer_0[1664] = in[210] | in[26]; 
    assign layer_0[1665] = in[25] | in[146]; 
    assign layer_0[1666] = in[149] & ~in[167]; 
    assign layer_0[1667] = ~in[58] | (in[58] & in[29]); 
    assign layer_0[1668] = in[186] & ~in[99]; 
    assign layer_0[1669] = ~(in[43] ^ in[75]); 
    assign layer_0[1670] = in[186] & ~in[198]; 
    assign layer_0[1671] = ~(in[243] ^ in[227]); 
    assign layer_0[1672] = ~(in[130] | in[131]); 
    assign layer_0[1673] = in[251] ^ in[204]; 
    assign layer_0[1674] = ~(in[37] ^ in[51]); 
    assign layer_0[1675] = ~(in[247] ^ in[137]); 
    assign layer_0[1676] = ~(in[246] ^ in[215]); 
    assign layer_0[1677] = ~in[55] | (in[102] & in[55]); 
    assign layer_0[1678] = in[90]; 
    assign layer_0[1679] = ~(in[159] | in[156]); 
    assign layer_0[1680] = in[199] ^ in[101]; 
    assign layer_0[1681] = ~(in[196] ^ in[38]); 
    assign layer_0[1682] = ~(in[115] ^ in[63]); 
    assign layer_0[1683] = ~(in[165] | in[199]); 
    assign layer_0[1684] = in[165] | in[179]; 
    assign layer_0[1685] = in[123] | in[203]; 
    assign layer_0[1686] = ~(in[147] | in[199]); 
    assign layer_0[1687] = ~(in[88] | in[94]); 
    assign layer_0[1688] = ~(in[131] ^ in[117]); 
    assign layer_0[1689] = ~(in[75] ^ in[27]); 
    assign layer_0[1690] = ~in[218] | (in[109] & in[218]); 
    assign layer_0[1691] = ~in[121]; 
    assign layer_0[1692] = ~(in[67] | in[72]); 
    assign layer_0[1693] = ~(in[221] ^ in[86]); 
    assign layer_0[1694] = in[137] & ~in[178]; 
    assign layer_0[1695] = in[231] | in[250]; 
    assign layer_0[1696] = in[221] ^ in[189]; 
    assign layer_0[1697] = ~(in[24] ^ in[126]); 
    assign layer_0[1698] = in[113] ^ in[100]; 
    assign layer_0[1699] = ~(in[109] | in[12]); 
    assign layer_0[1700] = in[133] ^ in[146]; 
    assign layer_0[1701] = in[145] | in[159]; 
    assign layer_0[1702] = ~(in[122] ^ in[166]); 
    assign layer_0[1703] = ~(in[236] | in[168]); 
    assign layer_0[1704] = ~(in[25] | in[143]); 
    assign layer_0[1705] = in[52] | in[83]; 
    assign layer_0[1706] = in[234] ^ in[219]; 
    assign layer_0[1707] = in[197] ^ in[53]; 
    assign layer_0[1708] = ~in[76] | (in[221] & in[76]); 
    assign layer_0[1709] = ~(in[186] ^ in[54]); 
    assign layer_0[1710] = ~(in[178] ^ in[165]); 
    assign layer_0[1711] = in[100] | in[72]; 
    assign layer_0[1712] = in[198] | in[213]; 
    assign layer_0[1713] = in[114] ^ in[101]; 
    assign layer_0[1714] = ~(in[220] ^ in[215]); 
    assign layer_0[1715] = ~in[196]; 
    assign layer_0[1716] = ~(in[162] | in[166]); 
    assign layer_0[1717] = ~(in[41] ^ in[243]); 
    assign layer_0[1718] = ~(in[117] | in[190]); 
    assign layer_0[1719] = in[108] ^ in[27]; 
    assign layer_0[1720] = ~in[219]; 
    assign layer_0[1721] = ~in[135] | (in[246] & in[135]); 
    assign layer_0[1722] = ~(in[154] | in[68]); 
    assign layer_0[1723] = ~(in[190] ^ in[126]); 
    assign layer_0[1724] = in[45] ^ in[230]; 
    assign layer_0[1725] = ~in[9]; 
    assign layer_0[1726] = in[243] | in[141]; 
    assign layer_0[1727] = ~(in[41] | in[72]); 
    assign layer_0[1728] = in[149] ^ in[147]; 
    assign layer_0[1729] = in[231] & ~in[184]; 
    assign layer_0[1730] = in[197] & ~in[22]; 
    assign layer_0[1731] = in[102]; 
    assign layer_0[1732] = ~(in[11] | in[251]); 
    assign layer_0[1733] = in[214] & ~in[85]; 
    assign layer_0[1734] = ~(in[88] ^ in[66]); 
    assign layer_0[1735] = ~(in[132] ^ in[103]); 
    assign layer_0[1736] = ~(in[232] | in[50]); 
    assign layer_0[1737] = ~(in[126] ^ in[108]); 
    assign layer_0[1738] = ~in[235]; 
    assign layer_0[1739] = in[182] ^ in[110]; 
    assign layer_0[1740] = ~in[136]; 
    assign layer_0[1741] = in[153] ^ in[122]; 
    assign layer_0[1742] = ~in[118]; 
    assign layer_0[1743] = in[134]; 
    assign layer_0[1744] = ~(in[165] | in[198]); 
    assign layer_0[1745] = in[232] ^ in[204]; 
    assign layer_0[1746] = ~in[216] | (in[146] & in[216]); 
    assign layer_0[1747] = in[125] ^ in[105]; 
    assign layer_0[1748] = ~(in[89] | in[172]); 
    assign layer_0[1749] = ~(in[140] ^ in[126]); 
    assign layer_0[1750] = in[230] ^ in[55]; 
    assign layer_0[1751] = ~(in[91] | in[170]); 
    assign layer_0[1752] = in[105] & ~in[54]; 
    assign layer_0[1753] = ~(in[63] | in[248]); 
    assign layer_0[1754] = in[228] | in[210]; 
    assign layer_0[1755] = in[129]; 
    assign layer_0[1756] = in[88] & ~in[108]; 
    assign layer_0[1757] = ~in[57] | (in[152] & in[57]); 
    assign layer_0[1758] = ~(in[213] ^ in[89]); 
    assign layer_0[1759] = ~in[38]; 
    assign layer_0[1760] = ~(in[211] | in[5]); 
    assign layer_0[1761] = in[147]; 
    assign layer_0[1762] = ~(in[174] ^ in[219]); 
    assign layer_0[1763] = ~(in[152] ^ in[47]); 
    assign layer_0[1764] = ~(in[243] ^ in[212]); 
    assign layer_0[1765] = ~(in[103] ^ in[139]); 
    assign layer_0[1766] = in[149] ^ in[102]; 
    assign layer_0[1767] = in[221] | in[194]; 
    assign layer_0[1768] = ~(in[43] ^ in[116]); 
    assign layer_0[1769] = ~(in[235] ^ in[203]); 
    assign layer_0[1770] = in[216] | in[22]; 
    assign layer_0[1771] = ~(in[73] ^ in[52]); 
    assign layer_0[1772] = ~(in[166] ^ in[198]); 
    assign layer_0[1773] = ~in[228]; 
    assign layer_0[1774] = in[216] ^ in[232]; 
    assign layer_0[1775] = in[121] | in[182]; 
    assign layer_0[1776] = in[104] ^ in[169]; 
    assign layer_0[1777] = in[180] | in[194]; 
    assign layer_0[1778] = in[196] & ~in[227]; 
    assign layer_0[1779] = in[21] ^ in[82]; 
    assign layer_0[1780] = in[11] | in[158]; 
    assign layer_0[1781] = in[183] & ~in[242]; 
    assign layer_0[1782] = in[24] ^ in[72]; 
    assign layer_0[1783] = in[55] & ~in[27]; 
    assign layer_0[1784] = in[230] | in[244]; 
    assign layer_0[1785] = ~(in[167] ^ in[119]); 
    assign layer_0[1786] = ~(in[130] | in[147]); 
    assign layer_0[1787] = ~(in[163] | in[90]); 
    assign layer_0[1788] = ~(in[190] ^ in[118]); 
    assign layer_0[1789] = ~(in[168] ^ in[150]); 
    assign layer_0[1790] = in[73] ^ in[42]; 
    assign layer_0[1791] = ~(in[77] ^ in[45]); 
    assign layer_0[1792] = in[47] | in[10]; 
    assign layer_0[1793] = in[233] | in[204]; 
    assign layer_0[1794] = ~(in[46] ^ in[93]); 
    assign layer_0[1795] = in[173] | in[75]; 
    assign layer_0[1796] = in[199] & ~in[85]; 
    assign layer_0[1797] = in[58] | in[90]; 
    assign layer_0[1798] = ~(in[119] ^ in[132]); 
    assign layer_0[1799] = in[73] ^ in[237]; 
    assign layer_0[1800] = ~(in[167] ^ in[211]); 
    assign layer_0[1801] = in[201] ^ in[182]; 
    assign layer_0[1802] = in[123] | in[140]; 
    assign layer_0[1803] = ~(in[172] | in[27]); 
    assign layer_0[1804] = in[35] ^ in[101]; 
    assign layer_0[1805] = ~in[42] | (in[219] & in[42]); 
    assign layer_0[1806] = in[46]; 
    assign layer_0[1807] = ~in[150] | (in[183] & in[150]); 
    assign layer_0[1808] = ~(in[60] ^ in[234]); 
    assign layer_0[1809] = in[151]; 
    assign layer_0[1810] = ~in[85]; 
    assign layer_0[1811] = ~(in[212] ^ in[82]); 
    assign layer_0[1812] = ~(in[149] ^ in[131]); 
    assign layer_0[1813] = in[34] | in[243]; 
    assign layer_0[1814] = ~in[137]; 
    assign layer_0[1815] = in[133] | in[69]; 
    assign layer_0[1816] = ~(in[147] ^ in[168]); 
    assign layer_0[1817] = in[140] ^ in[102]; 
    assign layer_0[1818] = in[83] ^ in[77]; 
    assign layer_0[1819] = ~(in[245] ^ in[217]); 
    assign layer_0[1820] = ~(in[205] ^ in[166]); 
    assign layer_0[1821] = ~(in[202] ^ in[248]); 
    assign layer_0[1822] = in[60] | in[104]; 
    assign layer_0[1823] = ~in[214] | (in[214] & in[105]); 
    assign layer_0[1824] = in[183] ^ in[214]; 
    assign layer_0[1825] = in[166] ^ in[201]; 
    assign layer_0[1826] = in[37] ^ in[198]; 
    assign layer_0[1827] = in[136] ^ in[22]; 
    assign layer_0[1828] = in[59] ^ in[183]; 
    assign layer_0[1829] = in[204] ^ in[173]; 
    assign layer_0[1830] = in[88] & ~in[106]; 
    assign layer_0[1831] = in[155] ^ in[182]; 
    assign layer_0[1832] = in[173] | in[204]; 
    assign layer_0[1833] = ~in[230] | (in[230] & in[183]); 
    assign layer_0[1834] = in[148] | in[130]; 
    assign layer_0[1835] = in[244] ^ in[34]; 
    assign layer_0[1836] = ~(in[41] ^ in[183]); 
    assign layer_0[1837] = in[197] ^ in[136]; 
    assign layer_0[1838] = ~in[149] | (in[149] & in[179]); 
    assign layer_0[1839] = in[36] | in[74]; 
    assign layer_0[1840] = in[100]; 
    assign layer_0[1841] = ~in[103]; 
    assign layer_0[1842] = ~(in[21] & in[213]); 
    assign layer_0[1843] = in[194] & ~in[81]; 
    assign layer_0[1844] = ~(in[235] ^ in[20]); 
    assign layer_0[1845] = ~(in[187] ^ in[205]); 
    assign layer_0[1846] = ~(in[107] ^ in[76]); 
    assign layer_0[1847] = in[90] & ~in[86]; 
    assign layer_0[1848] = in[61] ^ in[27]; 
    assign layer_0[1849] = in[131] & ~in[96]; 
    assign layer_0[1850] = in[11] ^ in[209]; 
    assign layer_0[1851] = ~in[152] | (in[152] & in[177]); 
    assign layer_0[1852] = in[251]; 
    assign layer_0[1853] = in[154] ^ in[135]; 
    assign layer_0[1854] = in[100] | in[156]; 
    assign layer_0[1855] = ~(in[245] | in[52]); 
    assign layer_0[1856] = in[47] | in[52]; 
    assign layer_0[1857] = ~(in[139] | in[156]); 
    assign layer_0[1858] = in[165] | in[120]; 
    assign layer_0[1859] = ~in[217] | (in[217] & in[39]); 
    assign layer_0[1860] = in[150] | in[27]; 
    assign layer_0[1861] = ~(in[184] & in[249]); 
    assign layer_0[1862] = in[251] ^ in[158]; 
    assign layer_0[1863] = in[93] & ~in[182]; 
    assign layer_0[1864] = in[196] ^ in[182]; 
    assign layer_0[1865] = ~(in[21] | in[138]); 
    assign layer_0[1866] = ~(in[68] ^ in[88]); 
    assign layer_0[1867] = ~in[165] | (in[123] & in[165]); 
    assign layer_0[1868] = in[41] & ~in[124]; 
    assign layer_0[1869] = in[84] ^ in[119]; 
    assign layer_0[1870] = ~(in[184] ^ in[138]); 
    assign layer_0[1871] = in[40] ^ in[87]; 
    assign layer_0[1872] = ~(in[61] ^ in[89]); 
    assign layer_0[1873] = ~(in[89] | in[243]); 
    assign layer_0[1874] = ~(in[228] ^ in[182]); 
    assign layer_0[1875] = in[107] ^ in[109]; 
    assign layer_0[1876] = ~in[229] | (in[180] & in[229]); 
    assign layer_0[1877] = ~(in[93] ^ in[105]); 
    assign layer_0[1878] = in[53]; 
    assign layer_0[1879] = ~(in[87] ^ in[42]); 
    assign layer_0[1880] = ~(in[177] | in[5]); 
    assign layer_0[1881] = ~(in[39] | in[39]); 
    assign layer_0[1882] = ~(in[74] ^ in[119]); 
    assign layer_0[1883] = in[165] & ~in[244]; 
    assign layer_0[1884] = in[198] | in[114]; 
    assign layer_0[1885] = in[167] ^ in[104]; 
    assign layer_0[1886] = ~(in[116] | in[113]); 
    assign layer_0[1887] = ~(in[201] ^ in[220]); 
    assign layer_0[1888] = ~(in[78] ^ in[56]); 
    assign layer_0[1889] = in[197] | in[198]; 
    assign layer_0[1890] = in[166] & ~in[85]; 
    assign layer_0[1891] = in[234] ^ in[219]; 
    assign layer_0[1892] = ~(in[22] | in[188]); 
    assign layer_0[1893] = ~(in[109] ^ in[120]); 
    assign layer_0[1894] = ~in[155] | (in[246] & in[155]); 
    assign layer_0[1895] = ~in[163] | (in[211] & in[163]); 
    assign layer_0[1896] = in[140] ^ in[157]; 
    assign layer_0[1897] = ~in[200] | (in[171] & in[200]); 
    assign layer_0[1898] = in[94] | in[76]; 
    assign layer_0[1899] = ~in[101] | (in[53] & in[101]); 
    assign layer_0[1900] = ~in[66]; 
    assign layer_0[1901] = in[5] ^ in[53]; 
    assign layer_0[1902] = in[245] & ~in[181]; 
    assign layer_0[1903] = in[69] & ~in[118]; 
    assign layer_0[1904] = in[198] ^ in[170]; 
    assign layer_0[1905] = in[118] ^ in[87]; 
    assign layer_0[1906] = ~(in[249] | in[221]); 
    assign layer_0[1907] = in[92] ^ in[189]; 
    assign layer_0[1908] = in[132]; 
    assign layer_0[1909] = in[242] | in[129]; 
    assign layer_0[1910] = in[165] ^ in[163]; 
    assign layer_0[1911] = ~(in[136] | in[168]); 
    assign layer_0[1912] = in[35] | in[181]; 
    assign layer_0[1913] = in[201] | in[232]; 
    assign layer_0[1914] = in[68] ^ in[230]; 
    assign layer_0[1915] = in[251]; 
    assign layer_0[1916] = in[210] | in[194]; 
    assign layer_0[1917] = ~in[234] | (in[135] & in[234]); 
    assign layer_0[1918] = in[90] | in[106]; 
    assign layer_0[1919] = ~(in[87] | in[72]); 
    assign layer_0[1920] = ~in[76] | (in[76] & in[165]); 
    assign layer_0[1921] = in[38] | in[205]; 
    assign layer_0[1922] = in[220] ^ in[9]; 
    assign layer_0[1923] = in[99] & ~in[78]; 
    assign layer_0[1924] = in[75]; 
    assign layer_0[1925] = ~(in[58] ^ in[11]); 
    assign layer_0[1926] = in[152] | in[121]; 
    assign layer_0[1927] = in[92] ^ in[73]; 
    assign layer_0[1928] = ~(in[38] ^ in[58]); 
    assign layer_0[1929] = ~in[53]; 
    assign layer_0[1930] = ~(in[116] ^ in[149]); 
    assign layer_0[1931] = ~(in[134] ^ in[248]); 
    assign layer_0[1932] = ~in[85] | (in[71] & in[85]); 
    assign layer_0[1933] = ~in[176]; 
    assign layer_0[1934] = in[89] | in[75]; 
    assign layer_0[1935] = in[180] | in[116]; 
    assign layer_0[1936] = in[92] ^ in[167]; 
    assign layer_0[1937] = ~(in[116] & in[84]); 
    assign layer_0[1938] = ~(in[129] | in[47]); 
    assign layer_0[1939] = in[175] | in[62]; 
    assign layer_0[1940] = in[171] & ~in[212]; 
    assign layer_0[1941] = ~(in[126] | in[116]); 
    assign layer_0[1942] = ~(in[27] ^ in[60]); 
    assign layer_0[1943] = in[177] ^ in[209]; 
    assign layer_0[1944] = ~(in[173] ^ in[242]); 
    assign layer_0[1945] = ~in[166] | (in[166] & in[212]); 
    assign layer_0[1946] = in[76] | in[123]; 
    assign layer_0[1947] = in[218] & ~in[98]; 
    assign layer_0[1948] = ~in[136] | (in[136] & in[202]); 
    assign layer_0[1949] = in[233] ^ in[212]; 
    assign layer_0[1950] = in[217] & ~in[210]; 
    assign layer_0[1951] = ~(in[225] | in[37]); 
    assign layer_0[1952] = in[241] ^ in[138]; 
    assign layer_0[1953] = in[73] ^ in[43]; 
    assign layer_0[1954] = ~(in[98] ^ in[88]); 
    assign layer_0[1955] = in[57] ^ in[25]; 
    assign layer_0[1956] = in[97] ^ in[98]; 
    assign layer_0[1957] = in[19]; 
    assign layer_0[1958] = in[22]; 
    assign layer_0[1959] = in[104] & ~in[186]; 
    assign layer_0[1960] = in[38] ^ in[70]; 
    assign layer_0[1961] = ~(in[141] | in[8]); 
    assign layer_0[1962] = in[176] | in[6]; 
    assign layer_0[1963] = ~(in[73] ^ in[235]); 
    assign layer_0[1964] = in[109] | in[70]; 
    assign layer_0[1965] = in[143]; 
    assign layer_0[1966] = in[166] ^ in[117]; 
    assign layer_0[1967] = in[163] ^ in[114]; 
    assign layer_0[1968] = ~(in[126] | in[195]); 
    assign layer_0[1969] = ~(in[167] & in[89]); 
    assign layer_0[1970] = ~(in[98] ^ in[85]); 
    assign layer_0[1971] = in[27] ^ in[57]; 
    assign layer_0[1972] = in[105] & ~in[72]; 
    assign layer_0[1973] = ~in[117] | (in[69] & in[117]); 
    assign layer_0[1974] = ~in[248] | (in[248] & in[153]); 
    assign layer_0[1975] = ~in[168] | (in[168] & in[163]); 
    assign layer_0[1976] = ~(in[201] ^ in[143]); 
    assign layer_0[1977] = in[103] ^ in[134]; 
    assign layer_0[1978] = ~(in[53] ^ in[99]); 
    assign layer_0[1979] = ~(in[119] ^ in[154]); 
    assign layer_0[1980] = in[78] | in[229]; 
    assign layer_0[1981] = ~(in[51] ^ in[37]); 
    assign layer_0[1982] = in[148] ^ in[28]; 
    assign layer_0[1983] = in[164] ^ in[199]; 
    assign layer_0[1984] = ~(in[99] | in[196]); 
    assign layer_0[1985] = in[75] | in[60]; 
    assign layer_0[1986] = in[141]; 
    assign layer_0[1987] = in[187] ^ in[196]; 
    assign layer_0[1988] = ~in[50] | (in[60] & in[50]); 
    assign layer_0[1989] = in[101]; 
    assign layer_0[1990] = in[214] | in[227]; 
    assign layer_0[1991] = ~(in[204] ^ in[201]); 
    assign layer_0[1992] = in[230]; 
    assign layer_0[1993] = in[173] | in[51]; 
    assign layer_0[1994] = in[152] & ~in[188]; 
    assign layer_0[1995] = in[191] | in[143]; 
    assign layer_0[1996] = in[203]; 
    assign layer_0[1997] = ~in[85] | (in[85] & in[120]); 
    assign layer_0[1998] = ~(in[173] ^ in[140]); 
    assign layer_0[1999] = in[197] | in[163]; 
    assign layer_0[2000] = in[107] ^ in[89]; 
    assign layer_0[2001] = ~(in[69] | in[199]); 
    assign layer_0[2002] = in[40] ^ in[177]; 
    assign layer_0[2003] = ~(in[84] | in[109]); 
    assign layer_0[2004] = in[177] & ~in[231]; 
    assign layer_0[2005] = in[212] & ~in[154]; 
    assign layer_0[2006] = in[231] | in[73]; 
    assign layer_0[2007] = ~(in[119] & in[54]); 
    assign layer_0[2008] = ~in[9] | (in[9] & in[173]); 
    assign layer_0[2009] = in[235]; 
    assign layer_0[2010] = in[6]; 
    assign layer_0[2011] = in[58] & ~in[54]; 
    assign layer_0[2012] = ~in[137] | (in[140] & in[137]); 
    assign layer_0[2013] = ~in[185]; 
    assign layer_0[2014] = in[86] & ~in[42]; 
    assign layer_0[2015] = in[212] ^ in[62]; 
    assign layer_0[2016] = ~in[133]; 
    assign layer_0[2017] = ~in[65]; 
    assign layer_0[2018] = ~(in[81] ^ in[34]); 
    assign layer_0[2019] = in[37] ^ in[101]; 
    assign layer_0[2020] = ~in[200] | (in[56] & in[200]); 
    assign layer_0[2021] = in[132] ^ in[118]; 
    assign layer_0[2022] = in[7] ^ in[20]; 
    assign layer_0[2023] = in[214] ^ in[166]; 
    assign layer_0[2024] = in[149] ^ in[146]; 
    assign layer_0[2025] = in[230] | in[228]; 
    assign layer_0[2026] = ~in[216] | (in[138] & in[216]); 
    assign layer_0[2027] = in[140] ^ in[109]; 
    assign layer_0[2028] = ~(in[200] & in[7]); 
    assign layer_0[2029] = in[88]; 
    assign layer_0[2030] = ~(in[247] | in[244]); 
    assign layer_0[2031] = ~(in[204] ^ in[22]); 
    assign layer_0[2032] = in[132] ^ in[165]; 
    assign layer_0[2033] = ~(in[94] ^ in[137]); 
    assign layer_0[2034] = ~in[152]; 
    assign layer_0[2035] = ~(in[181] | in[164]); 
    assign layer_0[2036] = ~(in[41] ^ in[72]); 
    assign layer_0[2037] = in[166] ^ in[201]; 
    assign layer_0[2038] = ~(in[197] ^ in[228]); 
    assign layer_0[2039] = in[146] ^ in[62]; 
    assign layer_0[2040] = ~(in[41] | in[120]); 
    assign layer_0[2041] = in[102] ^ in[117]; 
    assign layer_0[2042] = ~in[85] | (in[22] & in[85]); 
    assign layer_0[2043] = in[35] ^ in[235]; 
    assign layer_0[2044] = in[67] | in[106]; 
    assign layer_0[2045] = in[5] | in[162]; 
    assign layer_0[2046] = ~(in[45] | in[190]); 
    assign layer_0[2047] = ~(in[74] & in[26]); 
    assign layer_0[2048] = ~(in[215] | in[195]); 
    assign layer_0[2049] = in[183] | in[162]; 
    assign layer_0[2050] = ~(in[173] ^ in[118]); 
    assign layer_0[2051] = in[106] ^ in[179]; 
    assign layer_0[2052] = in[147] ^ in[118]; 
    assign layer_0[2053] = ~(in[123] ^ in[76]); 
    assign layer_0[2054] = ~in[118] | (in[118] & in[111]); 
    assign layer_0[2055] = ~(in[229] ^ in[214]); 
    assign layer_0[2056] = ~(in[184] ^ in[220]); 
    assign layer_0[2057] = in[205] | in[173]; 
    assign layer_0[2058] = in[103] | in[24]; 
    assign layer_0[2059] = in[187] ^ in[235]; 
    assign layer_0[2060] = in[41] ^ in[133]; 
    assign layer_0[2061] = in[166] ^ in[211]; 
    assign layer_0[2062] = in[204] | in[179]; 
    assign layer_0[2063] = in[5] | in[209]; 
    assign layer_0[2064] = in[118] ^ in[146]; 
    assign layer_0[2065] = in[194] ^ in[9]; 
    assign layer_0[2066] = ~(in[147] | in[63]); 
    assign layer_0[2067] = in[30] | in[212]; 
    assign layer_0[2068] = ~(in[103] ^ in[189]); 
    assign layer_0[2069] = ~(in[199] ^ in[133]); 
    assign layer_0[2070] = ~in[107]; 
    assign layer_0[2071] = in[141] ^ in[59]; 
    assign layer_0[2072] = ~(in[156] ^ in[250]); 
    assign layer_0[2073] = in[226] | in[37]; 
    assign layer_0[2074] = in[65]; 
    assign layer_0[2075] = in[200] ^ in[181]; 
    assign layer_0[2076] = in[116] ^ in[130]; 
    assign layer_0[2077] = in[142] | in[131]; 
    assign layer_0[2078] = in[188] | in[251]; 
    assign layer_0[2079] = in[57] ^ in[83]; 
    assign layer_0[2080] = ~(in[172] ^ in[118]); 
    assign layer_0[2081] = ~in[85] | (in[85] & in[193]); 
    assign layer_0[2082] = in[227] ^ in[243]; 
    assign layer_0[2083] = in[197] ^ in[71]; 
    assign layer_0[2084] = in[60] & in[247]; 
    assign layer_0[2085] = in[132] ^ in[40]; 
    assign layer_0[2086] = ~(in[52] ^ in[117]); 
    assign layer_0[2087] = ~in[180] | (in[180] & in[61]); 
    assign layer_0[2088] = ~(in[143] | in[141]); 
    assign layer_0[2089] = ~(in[76] ^ in[44]); 
    assign layer_0[2090] = ~in[103]; 
    assign layer_0[2091] = in[171]; 
    assign layer_0[2092] = ~(in[70] ^ in[84]); 
    assign layer_0[2093] = ~(in[196] ^ in[200]); 
    assign layer_0[2094] = ~(in[120] | in[136]); 
    assign layer_0[2095] = in[186] & ~in[86]; 
    assign layer_0[2096] = ~in[219] | (in[219] & in[181]); 
    assign layer_0[2097] = ~(in[202] | in[132]); 
    assign layer_0[2098] = ~in[189]; 
    assign layer_0[2099] = in[124] ^ in[183]; 
    assign layer_0[2100] = in[41] ^ in[73]; 
    assign layer_0[2101] = in[85] ^ in[181]; 
    assign layer_0[2102] = ~(in[206] ^ in[237]); 
    assign layer_0[2103] = in[59] & in[213]; 
    assign layer_0[2104] = ~(in[85] ^ in[70]); 
    assign layer_0[2105] = in[109] & ~in[79]; 
    assign layer_0[2106] = in[79] | in[248]; 
    assign layer_0[2107] = in[163] ^ in[181]; 
    assign layer_0[2108] = ~in[131] | (in[221] & in[131]); 
    assign layer_0[2109] = ~(in[202] ^ in[165]); 
    assign layer_0[2110] = in[150] ^ in[182]; 
    assign layer_0[2111] = ~in[233]; 
    assign layer_0[2112] = ~(in[168] ^ in[166]); 
    assign layer_0[2113] = in[122] & ~in[78]; 
    assign layer_0[2114] = in[74] & ~in[55]; 
    assign layer_0[2115] = in[38] & ~in[200]; 
    assign layer_0[2116] = ~in[135] | (in[241] & in[135]); 
    assign layer_0[2117] = ~(in[79] ^ in[221]); 
    assign layer_0[2118] = in[117] & ~in[141]; 
    assign layer_0[2119] = ~in[19]; 
    assign layer_0[2120] = in[77] | in[120]; 
    assign layer_0[2121] = ~in[41] | (in[41] & in[45]); 
    assign layer_0[2122] = ~(in[182] ^ in[164]); 
    assign layer_0[2123] = in[137] ^ in[182]; 
    assign layer_0[2124] = in[6] ^ in[221]; 
    assign layer_0[2125] = in[247] ^ in[150]; 
    assign layer_0[2126] = ~(in[185] ^ in[182]); 
    assign layer_0[2127] = ~in[86] | (in[234] & in[86]); 
    assign layer_0[2128] = ~(in[248] ^ in[219]); 
    assign layer_0[2129] = ~(in[166] ^ in[60]); 
    assign layer_0[2130] = ~in[200] | (in[71] & in[200]); 
    assign layer_0[2131] = ~in[140] | (in[140] & in[78]); 
    assign layer_0[2132] = ~(in[165] ^ in[150]); 
    assign layer_0[2133] = in[178] & ~in[109]; 
    assign layer_0[2134] = in[51] ^ in[197]; 
    assign layer_0[2135] = in[185] & ~in[66]; 
    assign layer_0[2136] = ~in[87] | (in[73] & in[87]); 
    assign layer_0[2137] = ~(in[24] ^ in[55]); 
    assign layer_0[2138] = in[50] ^ in[78]; 
    assign layer_0[2139] = in[74] ^ in[125]; 
    assign layer_0[2140] = in[71] ^ in[85]; 
    assign layer_0[2141] = ~(in[120] ^ in[134]); 
    assign layer_0[2142] = ~(in[70] | in[186]); 
    assign layer_0[2143] = ~(in[249] ^ in[235]); 
    assign layer_0[2144] = ~(in[105] ^ in[52]); 
    assign layer_0[2145] = in[27] ^ in[149]; 
    assign layer_0[2146] = ~in[26]; 
    assign layer_0[2147] = in[92] ^ in[89]; 
    assign layer_0[2148] = ~(in[194] | in[135]); 
    assign layer_0[2149] = in[98] | in[70]; 
    assign layer_0[2150] = ~(in[93] ^ in[167]); 
    assign layer_0[2151] = in[49] ^ in[46]; 
    assign layer_0[2152] = in[109] ^ in[111]; 
    assign layer_0[2153] = ~(in[86] | in[84]); 
    assign layer_0[2154] = ~(in[171] | in[203]); 
    assign layer_0[2155] = in[121] & ~in[140]; 
    assign layer_0[2156] = in[163] ^ in[165]; 
    assign layer_0[2157] = ~in[218]; 
    assign layer_0[2158] = in[54] | in[249]; 
    assign layer_0[2159] = in[23] & ~in[98]; 
    assign layer_0[2160] = ~in[197]; 
    assign layer_0[2161] = in[68] ^ in[82]; 
    assign layer_0[2162] = ~(in[199] ^ in[231]); 
    assign layer_0[2163] = in[26]; 
    assign layer_0[2164] = ~(in[166] ^ in[148]); 
    assign layer_0[2165] = ~(in[25] | in[42]); 
    assign layer_0[2166] = ~(in[156] | in[122]); 
    assign layer_0[2167] = ~(in[181] | in[20]); 
    assign layer_0[2168] = ~in[184] | (in[184] & in[243]); 
    assign layer_0[2169] = in[210] | in[215]; 
    assign layer_0[2170] = in[206] | in[28]; 
    assign layer_0[2171] = in[130]; 
    assign layer_0[2172] = ~(in[184] ^ in[99]); 
    assign layer_0[2173] = in[243] | in[97]; 
    assign layer_0[2174] = in[73] | in[97]; 
    assign layer_0[2175] = in[46] | in[29]; 
    assign layer_0[2176] = ~in[58] | (in[151] & in[58]); 
    assign layer_0[2177] = ~(in[22] | in[118]); 
    assign layer_0[2178] = ~(in[154] | in[156]); 
    assign layer_0[2179] = ~in[154]; 
    assign layer_0[2180] = in[37] ^ in[123]; 
    assign layer_0[2181] = in[23] & ~in[30]; 
    assign layer_0[2182] = ~(in[95] ^ in[93]); 
    assign layer_0[2183] = in[133] & ~in[250]; 
    assign layer_0[2184] = ~in[195]; 
    assign layer_0[2185] = in[218] | in[60]; 
    assign layer_0[2186] = ~in[139] | (in[139] & in[220]); 
    assign layer_0[2187] = in[119] | in[237]; 
    assign layer_0[2188] = in[200] ^ in[182]; 
    assign layer_0[2189] = in[10] | in[21]; 
    assign layer_0[2190] = ~in[131]; 
    assign layer_0[2191] = in[69] ^ in[22]; 
    assign layer_0[2192] = in[123]; 
    assign layer_0[2193] = in[133] ^ in[119]; 
    assign layer_0[2194] = in[178]; 
    assign layer_0[2195] = in[140] ^ in[105]; 
    assign layer_0[2196] = in[86]; 
    assign layer_0[2197] = in[138] | in[183]; 
    assign layer_0[2198] = in[251] | in[212]; 
    assign layer_0[2199] = ~in[151] | (in[107] & in[151]); 
    assign layer_0[2200] = ~(in[25] ^ in[158]); 
    assign layer_0[2201] = ~in[231]; 
    assign layer_0[2202] = ~in[186] | (in[122] & in[186]); 
    assign layer_0[2203] = in[6] ^ in[35]; 
    assign layer_0[2204] = in[162] | in[9]; 
    assign layer_0[2205] = in[136] ^ in[213]; 
    assign layer_0[2206] = ~in[154] | (in[154] & in[205]); 
    assign layer_0[2207] = ~(in[197] | in[196]); 
    assign layer_0[2208] = ~in[123] | (in[178] & in[123]); 
    assign layer_0[2209] = ~(in[163] | in[133]); 
    assign layer_0[2210] = ~(in[86] ^ in[90]); 
    assign layer_0[2211] = ~(in[85] ^ in[130]); 
    assign layer_0[2212] = in[115]; 
    assign layer_0[2213] = ~(in[119] ^ in[142]); 
    assign layer_0[2214] = ~(in[117] | in[163]); 
    assign layer_0[2215] = in[124] ^ in[70]; 
    assign layer_0[2216] = in[135] & in[167]; 
    assign layer_0[2217] = ~(in[45] | in[158]); 
    assign layer_0[2218] = in[76] & ~in[120]; 
    assign layer_0[2219] = ~(in[59] ^ in[103]); 
    assign layer_0[2220] = ~(in[134] | in[170]); 
    assign layer_0[2221] = in[192] | in[9]; 
    assign layer_0[2222] = in[142] ^ in[155]; 
    assign layer_0[2223] = ~(in[246] | in[193]); 
    assign layer_0[2224] = ~in[99] | (in[99] & in[197]); 
    assign layer_0[2225] = ~in[228] | (in[228] & in[69]); 
    assign layer_0[2226] = in[132] | in[146]; 
    assign layer_0[2227] = in[115]; 
    assign layer_0[2228] = in[137] | in[225]; 
    assign layer_0[2229] = in[103] & ~in[117]; 
    assign layer_0[2230] = ~(in[5] | in[137]); 
    assign layer_0[2231] = in[107] ^ in[137]; 
    assign layer_0[2232] = ~in[3] | (in[3] & in[119]); 
    assign layer_0[2233] = ~(in[217] | in[251]); 
    assign layer_0[2234] = ~(in[148] ^ in[196]); 
    assign layer_0[2235] = ~(in[217] | in[86]); 
    assign layer_0[2236] = in[53]; 
    assign layer_0[2237] = ~(in[153] ^ in[83]); 
    assign layer_0[2238] = in[212] ^ in[166]; 
    assign layer_0[2239] = in[59] | in[92]; 
    assign layer_0[2240] = ~in[57] | (in[131] & in[57]); 
    assign layer_0[2241] = ~(in[53] | in[229]); 
    assign layer_0[2242] = in[11] | in[251]; 
    assign layer_0[2243] = ~(in[168] ^ in[203]); 
    assign layer_0[2244] = in[121] ^ in[23]; 
    assign layer_0[2245] = in[155] & ~in[182]; 
    assign layer_0[2246] = in[9]; 
    assign layer_0[2247] = ~(in[212] | in[116]); 
    assign layer_0[2248] = in[67] | in[242]; 
    assign layer_0[2249] = in[138] ^ in[119]; 
    assign layer_0[2250] = in[198] ^ in[213]; 
    assign layer_0[2251] = in[120]; 
    assign layer_0[2252] = in[136]; 
    assign layer_0[2253] = in[249]; 
    assign layer_0[2254] = in[250] ^ in[168]; 
    assign layer_0[2255] = ~in[117] | (in[117] & in[75]); 
    assign layer_0[2256] = in[187] ^ in[136]; 
    assign layer_0[2257] = ~(in[236] | in[203]); 
    assign layer_0[2258] = ~in[189] | (in[189] & in[157]); 
    assign layer_0[2259] = in[145]; 
    assign layer_0[2260] = in[189] | in[204]; 
    assign layer_0[2261] = ~in[169]; 
    assign layer_0[2262] = ~(in[197] ^ in[247]); 
    assign layer_0[2263] = in[83] | in[65]; 
    assign layer_0[2264] = ~(in[175] | in[5]); 
    assign layer_0[2265] = ~in[218] | (in[183] & in[218]); 
    assign layer_0[2266] = in[90] & ~in[116]; 
    assign layer_0[2267] = ~(in[106] ^ in[137]); 
    assign layer_0[2268] = in[252] | in[184]; 
    assign layer_0[2269] = ~(in[100] ^ in[98]); 
    assign layer_0[2270] = in[88] & ~in[41]; 
    assign layer_0[2271] = ~(in[242] | in[5]); 
    assign layer_0[2272] = ~(in[57] ^ in[59]); 
    assign layer_0[2273] = ~(in[116] | in[101]); 
    assign layer_0[2274] = ~(in[123] ^ in[137]); 
    assign layer_0[2275] = ~(in[55] | in[118]); 
    assign layer_0[2276] = in[136] ^ in[104]; 
    assign layer_0[2277] = ~(in[245] | in[166]); 
    assign layer_0[2278] = in[77] & ~in[137]; 
    assign layer_0[2279] = ~(in[95] ^ in[61]); 
    assign layer_0[2280] = ~(in[134] & in[163]); 
    assign layer_0[2281] = ~(in[249] ^ in[218]); 
    assign layer_0[2282] = ~in[136] | (in[44] & in[136]); 
    assign layer_0[2283] = ~(in[243] ^ in[129]); 
    assign layer_0[2284] = ~in[170] | (in[219] & in[170]); 
    assign layer_0[2285] = ~(in[117] ^ in[134]); 
    assign layer_0[2286] = in[36] ^ in[117]; 
    assign layer_0[2287] = ~(in[135] ^ in[140]); 
    assign layer_0[2288] = in[167] ^ in[198]; 
    assign layer_0[2289] = in[106] | in[170]; 
    assign layer_0[2290] = ~(in[114] | in[244]); 
    assign layer_0[2291] = ~(in[185] ^ in[232]); 
    assign layer_0[2292] = ~(in[155] | in[123]); 
    assign layer_0[2293] = ~(in[22] ^ in[136]); 
    assign layer_0[2294] = in[177] | in[65]; 
    assign layer_0[2295] = ~(in[201] | in[186]); 
    assign layer_0[2296] = ~in[215] | (in[245] & in[215]); 
    assign layer_0[2297] = in[57]; 
    assign layer_0[2298] = in[22] | in[221]; 
    assign layer_0[2299] = in[170] ^ in[156]; 
    assign layer_0[2300] = in[156] ^ in[122]; 
    assign layer_0[2301] = ~(in[181] | in[164]); 
    assign layer_0[2302] = ~(in[26] ^ in[193]); 
    assign layer_0[2303] = ~in[137] | (in[137] & in[130]); 
    assign layer_0[2304] = in[146] ^ in[148]; 
    assign layer_0[2305] = ~(in[166] ^ in[244]); 
    assign layer_0[2306] = ~(in[156] | in[98]); 
    assign layer_0[2307] = ~(in[29] | in[184]); 
    assign layer_0[2308] = in[101] & in[214]; 
    assign layer_0[2309] = in[108] & ~in[214]; 
    assign layer_0[2310] = in[114]; 
    assign layer_0[2311] = in[142] | in[137]; 
    assign layer_0[2312] = in[219] | in[243]; 
    assign layer_0[2313] = ~(in[148] | in[146]); 
    assign layer_0[2314] = ~(in[196] | in[198]); 
    assign layer_0[2315] = ~(in[251] ^ in[137]); 
    assign layer_0[2316] = in[101] & ~in[56]; 
    assign layer_0[2317] = ~(in[34] ^ in[65]); 
    assign layer_0[2318] = ~(in[41] ^ in[82]); 
    assign layer_0[2319] = ~in[217] | (in[106] & in[217]); 
    assign layer_0[2320] = in[219] ^ in[251]; 
    assign layer_0[2321] = ~(in[196] | in[188]); 
    assign layer_0[2322] = ~(in[219] & in[137]); 
    assign layer_0[2323] = in[211] ^ in[106]; 
    assign layer_0[2324] = ~in[233] | (in[230] & in[233]); 
    assign layer_0[2325] = in[223] | in[79]; 
    assign layer_0[2326] = in[83] | in[177]; 
    assign layer_0[2327] = ~(in[217] ^ in[232]); 
    assign layer_0[2328] = in[66] ^ in[93]; 
    assign layer_0[2329] = in[26] | in[162]; 
    assign layer_0[2330] = ~(in[106] | in[19]); 
    assign layer_0[2331] = in[53]; 
    assign layer_0[2332] = ~in[217] | (in[217] & in[72]); 
    assign layer_0[2333] = in[77]; 
    assign layer_0[2334] = in[69] ^ in[102]; 
    assign layer_0[2335] = ~(in[166] | in[151]); 
    assign layer_0[2336] = ~(in[115] ^ in[100]); 
    assign layer_0[2337] = ~(in[155] | in[53]); 
    assign layer_0[2338] = in[56]; 
    assign layer_0[2339] = ~(in[182] & in[150]); 
    assign layer_0[2340] = in[154] ^ in[12]; 
    assign layer_0[2341] = in[125]; 
    assign layer_0[2342] = in[177] | in[25]; 
    assign layer_0[2343] = ~(in[41] ^ in[113]); 
    assign layer_0[2344] = ~(in[28] ^ in[26]); 
    assign layer_0[2345] = in[190] | in[205]; 
    assign layer_0[2346] = in[211] | in[180]; 
    assign layer_0[2347] = in[120] & ~in[37]; 
    assign layer_0[2348] = ~(in[111] | in[142]); 
    assign layer_0[2349] = in[152] | in[221]; 
    assign layer_0[2350] = ~(in[121] | in[154]); 
    assign layer_0[2351] = in[124] & in[43]; 
    assign layer_0[2352] = ~in[74]; 
    assign layer_0[2353] = ~(in[28] | in[8]); 
    assign layer_0[2354] = in[74] ^ in[72]; 
    assign layer_0[2355] = ~(in[70] ^ in[100]); 
    assign layer_0[2356] = ~in[152] | (in[252] & in[152]); 
    assign layer_0[2357] = in[177] | in[88]; 
    assign layer_0[2358] = in[41] ^ in[57]; 
    assign layer_0[2359] = in[45] | in[65]; 
    assign layer_0[2360] = ~(in[54] | in[93]); 
    assign layer_0[2361] = ~(in[124] | in[91]); 
    assign layer_0[2362] = in[118]; 
    assign layer_0[2363] = ~(in[102] ^ in[117]); 
    assign layer_0[2364] = in[88] ^ in[57]; 
    assign layer_0[2365] = in[121] ^ in[166]; 
    assign layer_0[2366] = in[70] ^ in[74]; 
    assign layer_0[2367] = in[28] ^ in[73]; 
    assign layer_0[2368] = in[39] & ~in[118]; 
    assign layer_0[2369] = in[27] | in[179]; 
    assign layer_0[2370] = ~(in[157] ^ in[102]); 
    assign layer_0[2371] = in[67] | in[156]; 
    assign layer_0[2372] = in[171] ^ in[140]; 
    assign layer_0[2373] = ~(in[193] ^ in[190]); 
    assign layer_0[2374] = ~(in[244] ^ in[247]); 
    assign layer_0[2375] = in[225] | in[187]; 
    assign layer_0[2376] = in[148] ^ in[90]; 
    assign layer_0[2377] = in[156]; 
    assign layer_0[2378] = in[95] ^ in[39]; 
    assign layer_0[2379] = in[57] ^ in[27]; 
    assign layer_0[2380] = in[76] | in[168]; 
    assign layer_0[2381] = ~(in[183] | in[120]); 
    assign layer_0[2382] = ~in[40] | (in[40] & in[10]); 
    assign layer_0[2383] = ~(in[179] ^ in[205]); 
    assign layer_0[2384] = ~in[228]; 
    assign layer_0[2385] = ~(in[53] ^ in[21]); 
    assign layer_0[2386] = ~(in[234] & in[54]); 
    assign layer_0[2387] = ~(in[101] | in[37]); 
    assign layer_0[2388] = ~(in[94] ^ in[165]); 
    assign layer_0[2389] = in[137] | in[139]; 
    assign layer_0[2390] = in[185] ^ in[119]; 
    assign layer_0[2391] = ~(in[94] | in[183]); 
    assign layer_0[2392] = ~(in[140] & in[125]); 
    assign layer_0[2393] = ~(in[40] | in[55]); 
    assign layer_0[2394] = in[181] ^ in[211]; 
    assign layer_0[2395] = ~in[123]; 
    assign layer_0[2396] = in[172] ^ in[50]; 
    assign layer_0[2397] = ~(in[187] | in[20]); 
    assign layer_0[2398] = in[86] & ~in[206]; 
    assign layer_0[2399] = in[120] & in[139]; 
    assign layer_0[2400] = in[145]; 
    assign layer_0[2401] = in[210] & ~in[92]; 
    assign layer_0[2402] = ~in[168]; 
    assign layer_0[2403] = in[163] ^ in[165]; 
    assign layer_0[2404] = in[155] ^ in[252]; 
    assign layer_0[2405] = in[90] ^ in[189]; 
    assign layer_0[2406] = ~in[143]; 
    assign layer_0[2407] = ~(in[131] ^ in[177]); 
    assign layer_0[2408] = in[104] | in[119]; 
    assign layer_0[2409] = ~in[122] | (in[122] & in[172]); 
    assign layer_0[2410] = in[116] ^ in[213]; 
    assign layer_0[2411] = in[121] ^ in[183]; 
    assign layer_0[2412] = in[184] ^ in[44]; 
    assign layer_0[2413] = ~(in[170] ^ in[195]); 
    assign layer_0[2414] = ~(in[119] | in[134]); 
    assign layer_0[2415] = ~(in[170] ^ in[93]); 
    assign layer_0[2416] = in[116] | in[22]; 
    assign layer_0[2417] = in[230] ^ in[244]; 
    assign layer_0[2418] = ~(in[89] ^ in[53]); 
    assign layer_0[2419] = ~(in[198] ^ in[30]); 
    assign layer_0[2420] = in[178] | in[28]; 
    assign layer_0[2421] = ~(in[74] ^ in[172]); 
    assign layer_0[2422] = in[21] ^ in[24]; 
    assign layer_0[2423] = in[41] & in[55]; 
    assign layer_0[2424] = in[89] ^ in[91]; 
    assign layer_0[2425] = in[37] | in[24]; 
    assign layer_0[2426] = ~(in[236] ^ in[146]); 
    assign layer_0[2427] = ~(in[220] ^ in[173]); 
    assign layer_0[2428] = ~(in[167] | in[151]); 
    assign layer_0[2429] = in[228] ^ in[177]; 
    assign layer_0[2430] = ~in[245] | (in[165] & in[245]); 
    assign layer_0[2431] = in[245] & ~in[55]; 
    assign layer_0[2432] = in[153] & ~in[53]; 
    assign layer_0[2433] = ~(in[78] | in[98]); 
    assign layer_0[2434] = ~(in[197] ^ in[179]); 
    assign layer_0[2435] = ~(in[7] | in[210]); 
    assign layer_0[2436] = in[58] ^ in[89]; 
    assign layer_0[2437] = ~(in[150] ^ in[152]); 
    assign layer_0[2438] = ~(in[93] ^ in[151]); 
    assign layer_0[2439] = in[92] & ~in[151]; 
    assign layer_0[2440] = in[38] ^ in[104]; 
    assign layer_0[2441] = ~in[57]; 
    assign layer_0[2442] = ~(in[122] ^ in[197]); 
    assign layer_0[2443] = ~(in[154] ^ in[119]); 
    assign layer_0[2444] = in[67]; 
    assign layer_0[2445] = ~(in[246] ^ in[214]); 
    assign layer_0[2446] = ~(in[165] | in[99]); 
    assign layer_0[2447] = in[219]; 
    assign layer_0[2448] = ~(in[42] | in[52]); 
    assign layer_0[2449] = in[90] ^ in[94]; 
    assign layer_0[2450] = in[235] ^ in[206]; 
    assign layer_0[2451] = in[142] & in[57]; 
    assign layer_0[2452] = ~(in[79] | in[235]); 
    assign layer_0[2453] = in[106] ^ in[73]; 
    assign layer_0[2454] = ~(in[108] & in[75]); 
    assign layer_0[2455] = ~(in[131] | in[43]); 
    assign layer_0[2456] = ~in[230] | (in[245] & in[230]); 
    assign layer_0[2457] = in[92] ^ in[94]; 
    assign layer_0[2458] = ~(in[63] | in[130]); 
    assign layer_0[2459] = ~(in[157] | in[185]); 
    assign layer_0[2460] = in[202] ^ in[234]; 
    assign layer_0[2461] = in[40] ^ in[164]; 
    assign layer_0[2462] = in[118] ^ in[83]; 
    assign layer_0[2463] = in[135] ^ in[85]; 
    assign layer_0[2464] = in[150] | in[131]; 
    assign layer_0[2465] = in[183] ^ in[155]; 
    assign layer_0[2466] = ~(in[201] ^ in[84]); 
    assign layer_0[2467] = in[87] & ~in[131]; 
    assign layer_0[2468] = ~(in[86] | in[113]); 
    assign layer_0[2469] = ~in[168] | (in[229] & in[168]); 
    assign layer_0[2470] = ~in[5]; 
    assign layer_0[2471] = in[100] | in[78]; 
    assign layer_0[2472] = in[146] | in[164]; 
    assign layer_0[2473] = in[114] | in[153]; 
    assign layer_0[2474] = ~(in[77] ^ in[78]); 
    assign layer_0[2475] = ~(in[143] | in[74]); 
    assign layer_0[2476] = in[211]; 
    assign layer_0[2477] = ~in[86]; 
    assign layer_0[2478] = in[182]; 
    assign layer_0[2479] = ~(in[194] ^ in[197]); 
    assign layer_0[2480] = in[119] | in[141]; 
    assign layer_0[2481] = ~in[137] | (in[137] & in[193]); 
    assign layer_0[2482] = ~(in[120] ^ in[232]); 
    assign layer_0[2483] = in[46] ^ in[243]; 
    assign layer_0[2484] = ~(in[113] ^ in[73]); 
    assign layer_0[2485] = in[42] ^ in[73]; 
    assign layer_0[2486] = in[226] ^ in[72]; 
    assign layer_0[2487] = ~(in[6] | in[19]); 
    assign layer_0[2488] = in[42] ^ in[68]; 
    assign layer_0[2489] = ~(in[212] ^ in[198]); 
    assign layer_0[2490] = ~in[164]; 
    assign layer_0[2491] = ~in[105] | (in[150] & in[105]); 
    assign layer_0[2492] = in[183] & ~in[210]; 
    assign layer_0[2493] = in[103] | in[165]; 
    assign layer_0[2494] = in[251]; 
    assign layer_0[2495] = in[108] ^ in[215]; 
    assign layer_0[2496] = ~(in[8] | in[148]); 
    assign layer_0[2497] = in[213] & ~in[60]; 
    assign layer_0[2498] = in[165] | in[148]; 
    assign layer_0[2499] = ~(in[27] & in[87]); 
    assign layer_0[2500] = in[175] ^ in[194]; 
    assign layer_0[2501] = ~in[182] | (in[182] & in[103]); 
    assign layer_0[2502] = ~(in[133] | in[204]); 
    assign layer_0[2503] = in[213] ^ in[5]; 
    assign layer_0[2504] = ~in[203] | (in[80] & in[203]); 
    assign layer_0[2505] = in[152]; 
    assign layer_0[2506] = ~(in[35] ^ in[185]); 
    assign layer_0[2507] = ~in[103] | (in[103] & in[189]); 
    assign layer_0[2508] = ~(in[156] ^ in[68]); 
    assign layer_0[2509] = ~(in[145] | in[242]); 
    assign layer_0[2510] = ~(in[204] | in[52]); 
    assign layer_0[2511] = ~(in[100] ^ in[86]); 
    assign layer_0[2512] = ~(in[164] | in[143]); 
    assign layer_0[2513] = ~(in[246] ^ in[211]); 
    assign layer_0[2514] = ~(in[190] | in[175]); 
    assign layer_0[2515] = ~in[206]; 
    assign layer_0[2516] = ~(in[158] | in[171]); 
    assign layer_0[2517] = ~in[104] | (in[104] & in[148]); 
    assign layer_0[2518] = in[197] ^ in[138]; 
    assign layer_0[2519] = ~(in[134] | in[75]); 
    assign layer_0[2520] = ~(in[189] ^ in[133]); 
    assign layer_0[2521] = ~in[171] | (in[134] & in[171]); 
    assign layer_0[2522] = ~(in[9] | in[68]); 
    assign layer_0[2523] = ~(in[63] ^ in[46]); 
    assign layer_0[2524] = ~(in[249] ^ in[235]); 
    assign layer_0[2525] = in[52] ^ in[83]; 
    assign layer_0[2526] = ~in[151] | (in[151] & in[214]); 
    assign layer_0[2527] = ~(in[141] ^ in[59]); 
    assign layer_0[2528] = in[231] ^ in[200]; 
    assign layer_0[2529] = ~in[118] | (in[118] & in[91]); 
    assign layer_0[2530] = in[105] & ~in[222]; 
    assign layer_0[2531] = in[229] | in[247]; 
    assign layer_0[2532] = ~in[215] | (in[215] & in[131]); 
    assign layer_0[2533] = in[116] | in[159]; 
    assign layer_0[2534] = in[188] ^ in[89]; 
    assign layer_0[2535] = in[116] | in[87]; 
    assign layer_0[2536] = in[59] | in[92]; 
    assign layer_0[2537] = ~(in[185] | in[115]); 
    assign layer_0[2538] = ~(in[198] ^ in[140]); 
    assign layer_0[2539] = ~in[137] | (in[213] & in[137]); 
    assign layer_0[2540] = in[150] | in[37]; 
    assign layer_0[2541] = ~in[84] | (in[102] & in[84]); 
    assign layer_0[2542] = in[162] | in[164]; 
    assign layer_0[2543] = in[8]; 
    assign layer_0[2544] = ~(in[196] ^ in[158]); 
    assign layer_0[2545] = in[91] ^ in[60]; 
    assign layer_0[2546] = ~(in[49] | in[71]); 
    assign layer_0[2547] = in[210] ^ in[165]; 
    assign layer_0[2548] = in[137] ^ in[105]; 
    assign layer_0[2549] = in[249] ^ in[131]; 
    assign layer_0[2550] = in[189] ^ in[170]; 
    assign layer_0[2551] = in[166] ^ in[119]; 
    assign layer_0[2552] = ~(in[101] ^ in[114]); 
    assign layer_0[2553] = in[118]; 
    assign layer_0[2554] = in[53] ^ in[200]; 
    assign layer_0[2555] = ~in[72] | (in[180] & in[72]); 
    assign layer_0[2556] = in[117]; 
    assign layer_0[2557] = in[55] & ~in[85]; 
    assign layer_0[2558] = in[172] ^ in[74]; 
    assign layer_0[2559] = in[39] ^ in[8]; 
    assign layer_0[2560] = in[94] & in[117]; 
    assign layer_0[2561] = in[119] | in[195]; 
    assign layer_0[2562] = in[78] | in[26]; 
    assign layer_0[2563] = ~(in[213] | in[53]); 
    assign layer_0[2564] = in[118] ^ in[204]; 
    assign layer_0[2565] = in[87] | in[98]; 
    assign layer_0[2566] = ~in[185] | (in[218] & in[185]); 
    assign layer_0[2567] = in[90] ^ in[138]; 
    assign layer_0[2568] = in[24] | in[92]; 
    assign layer_0[2569] = in[169] ^ in[195]; 
    assign layer_0[2570] = ~(in[116] | in[108]); 
    assign layer_0[2571] = in[246] | in[227]; 
    assign layer_0[2572] = ~(in[94] | in[242]); 
    assign layer_0[2573] = in[136] | in[35]; 
    assign layer_0[2574] = in[251] ^ in[151]; 
    assign layer_0[2575] = ~(in[105] ^ in[168]); 
    assign layer_0[2576] = ~(in[171] ^ in[108]); 
    assign layer_0[2577] = ~(in[53] ^ in[92]); 
    assign layer_0[2578] = in[59] & ~in[26]; 
    assign layer_0[2579] = in[38] ^ in[54]; 
    assign layer_0[2580] = ~in[247] | (in[247] & in[213]); 
    assign layer_0[2581] = ~(in[72] ^ in[74]); 
    assign layer_0[2582] = in[119] ^ in[71]; 
    assign layer_0[2583] = ~(in[78] ^ in[76]); 
    assign layer_0[2584] = ~in[36] | (in[36] & in[74]); 
    assign layer_0[2585] = in[166] | in[115]; 
    assign layer_0[2586] = in[65] ^ in[94]; 
    assign layer_0[2587] = ~(in[136] ^ in[140]); 
    assign layer_0[2588] = ~in[242]; 
    assign layer_0[2589] = ~(in[103] ^ in[171]); 
    assign layer_0[2590] = in[132] ^ in[115]; 
    assign layer_0[2591] = ~(in[103] | in[205]); 
    assign layer_0[2592] = in[168] & ~in[229]; 
    assign layer_0[2593] = in[27] ^ in[61]; 
    assign layer_0[2594] = in[153]; 
    assign layer_0[2595] = ~(in[227] ^ in[51]); 
    assign layer_0[2596] = in[142] | in[236]; 
    assign layer_0[2597] = in[150] ^ in[152]; 
    assign layer_0[2598] = ~(in[106] ^ in[137]); 
    assign layer_0[2599] = ~(in[151] ^ in[217]); 
    assign layer_0[2600] = in[101] & ~in[53]; 
    assign layer_0[2601] = ~(in[123] | in[44]); 
    assign layer_0[2602] = ~in[63] | (in[63] & in[140]); 
    assign layer_0[2603] = in[103] & ~in[34]; 
    assign layer_0[2604] = ~(in[74] ^ in[106]); 
    assign layer_0[2605] = in[140] & ~in[186]; 
    assign layer_0[2606] = ~(in[242] | in[156]); 
    assign layer_0[2607] = ~(in[214] & in[232]); 
    assign layer_0[2608] = in[249] ^ in[60]; 
    assign layer_0[2609] = in[168]; 
    assign layer_0[2610] = in[179] | in[203]; 
    assign layer_0[2611] = in[58] ^ in[26]; 
    assign layer_0[2612] = in[148] ^ in[170]; 
    assign layer_0[2613] = in[71] ^ in[120]; 
    assign layer_0[2614] = ~(in[196] ^ in[131]); 
    assign layer_0[2615] = ~(in[147] ^ in[130]); 
    assign layer_0[2616] = in[221] | in[27]; 
    assign layer_0[2617] = ~in[145]; 
    assign layer_0[2618] = in[103] & in[73]; 
    assign layer_0[2619] = ~(in[86] | in[54]); 
    assign layer_0[2620] = ~(in[217] | in[187]); 
    assign layer_0[2621] = ~(in[195] | in[68]); 
    assign layer_0[2622] = ~in[229]; 
    assign layer_0[2623] = in[138] & ~in[164]; 
    assign layer_0[2624] = ~in[185] | (in[162] & in[185]); 
    assign layer_0[2625] = ~(in[138] ^ in[121]); 
    assign layer_0[2626] = ~(in[228] ^ in[198]); 
    assign layer_0[2627] = in[42] ^ in[89]; 
    assign layer_0[2628] = ~in[200] | (in[200] & in[42]); 
    assign layer_0[2629] = in[56] ^ in[219]; 
    assign layer_0[2630] = in[190] & ~in[73]; 
    assign layer_0[2631] = in[131] | in[226]; 
    assign layer_0[2632] = ~in[232]; 
    assign layer_0[2633] = in[103] ^ in[117]; 
    assign layer_0[2634] = ~in[179] | (in[179] & in[150]); 
    assign layer_0[2635] = ~(in[195] ^ in[248]); 
    assign layer_0[2636] = ~(in[87] ^ in[101]); 
    assign layer_0[2637] = in[56] ^ in[87]; 
    assign layer_0[2638] = ~(in[100] | in[41]); 
    assign layer_0[2639] = ~in[19]; 
    assign layer_0[2640] = in[182] ^ in[180]; 
    assign layer_0[2641] = in[40] | in[118]; 
    assign layer_0[2642] = ~(in[241] | in[142]); 
    assign layer_0[2643] = ~in[148] | (in[148] & in[183]); 
    assign layer_0[2644] = in[186]; 
    assign layer_0[2645] = in[151] ^ in[180]; 
    assign layer_0[2646] = in[210] | in[111]; 
    assign layer_0[2647] = in[71] | in[79]; 
    assign layer_0[2648] = in[86] | in[65]; 
    assign layer_0[2649] = ~(in[173] ^ in[204]); 
    assign layer_0[2650] = in[149] ^ in[103]; 
    assign layer_0[2651] = in[73] & ~in[151]; 
    assign layer_0[2652] = in[115] ^ in[101]; 
    assign layer_0[2653] = in[105] ^ in[92]; 
    assign layer_0[2654] = ~(in[180] ^ in[198]); 
    assign layer_0[2655] = in[177] ^ in[166]; 
    assign layer_0[2656] = ~(in[230] ^ in[215]); 
    assign layer_0[2657] = in[221] ^ in[179]; 
    assign layer_0[2658] = in[107] ^ in[139]; 
    assign layer_0[2659] = in[213] | in[198]; 
    assign layer_0[2660] = ~(in[123] ^ in[121]); 
    assign layer_0[2661] = in[143]; 
    assign layer_0[2662] = in[177] ^ in[7]; 
    assign layer_0[2663] = ~(in[26] ^ in[73]); 
    assign layer_0[2664] = ~in[233]; 
    assign layer_0[2665] = ~in[85] | (in[85] & in[200]); 
    assign layer_0[2666] = in[116] ^ in[114]; 
    assign layer_0[2667] = in[70] | in[45]; 
    assign layer_0[2668] = ~(in[36] | in[47]); 
    assign layer_0[2669] = in[132] | in[202]; 
    assign layer_0[2670] = in[76] ^ in[182]; 
    assign layer_0[2671] = in[247] & ~in[92]; 
    assign layer_0[2672] = ~(in[74] ^ in[72]); 
    assign layer_0[2673] = ~(in[149] | in[132]); 
    assign layer_0[2674] = ~in[137] | (in[30] & in[137]); 
    assign layer_0[2675] = in[137] ^ in[121]; 
    assign layer_0[2676] = 1'b0; 
    assign layer_0[2677] = in[91] & ~in[211]; 
    assign layer_0[2678] = ~(in[209] ^ in[156]); 
    assign layer_0[2679] = ~(in[228] | in[39]); 
    assign layer_0[2680] = ~in[42] | (in[181] & in[42]); 
    assign layer_0[2681] = ~(in[59] ^ in[93]); 
    assign layer_0[2682] = in[88] ^ in[175]; 
    assign layer_0[2683] = in[149]; 
    assign layer_0[2684] = in[119] ^ in[133]; 
    assign layer_0[2685] = ~(in[46] ^ in[29]); 
    assign layer_0[2686] = in[218] ^ in[182]; 
    assign layer_0[2687] = in[216] & ~in[67]; 
    assign layer_0[2688] = ~in[143] | (in[235] & in[143]); 
    assign layer_0[2689] = in[45] ^ in[70]; 
    assign layer_0[2690] = in[119] ^ in[132]; 
    assign layer_0[2691] = ~(in[76] ^ in[74]); 
    assign layer_0[2692] = ~(in[124] ^ in[157]); 
    assign layer_0[2693] = ~in[142] | (in[138] & in[142]); 
    assign layer_0[2694] = in[134] ^ in[164]; 
    assign layer_0[2695] = ~in[72] | (in[167] & in[72]); 
    assign layer_0[2696] = in[131] | in[130]; 
    assign layer_0[2697] = ~(in[148] ^ in[167]); 
    assign layer_0[2698] = ~in[90] | (in[90] & in[119]); 
    assign layer_0[2699] = ~in[110]; 
    assign layer_0[2700] = ~in[193]; 
    assign layer_0[2701] = in[236] | in[249]; 
    assign layer_0[2702] = in[149] | in[151]; 
    assign layer_0[2703] = in[199] | in[85]; 
    assign layer_0[2704] = in[57] & ~in[121]; 
    assign layer_0[2705] = ~in[37]; 
    assign layer_0[2706] = ~in[131] | (in[148] & in[131]); 
    assign layer_0[2707] = in[70] ^ in[23]; 
    assign layer_0[2708] = ~(in[77] | in[72]); 
    assign layer_0[2709] = in[102] & ~in[235]; 
    assign layer_0[2710] = in[149] ^ in[181]; 
    assign layer_0[2711] = ~in[135] | (in[8] & in[135]); 
    assign layer_0[2712] = ~(in[23] ^ in[106]); 
    assign layer_0[2713] = ~(in[75] | in[90]); 
    assign layer_0[2714] = in[84]; 
    assign layer_0[2715] = ~(in[210] | in[227]); 
    assign layer_0[2716] = in[27] ^ in[26]; 
    assign layer_0[2717] = in[141] ^ in[102]; 
    assign layer_0[2718] = in[181] | in[109]; 
    assign layer_0[2719] = in[101] & ~in[191]; 
    assign layer_0[2720] = in[150] & ~in[155]; 
    assign layer_0[2721] = in[196] ^ in[203]; 
    assign layer_0[2722] = in[107] | in[44]; 
    assign layer_0[2723] = in[122] ^ in[155]; 
    assign layer_0[2724] = in[97] & ~in[201]; 
    assign layer_0[2725] = in[77] ^ in[88]; 
    assign layer_0[2726] = ~(in[197] | in[195]); 
    assign layer_0[2727] = in[194] ^ in[212]; 
    assign layer_0[2728] = ~(in[199] ^ in[201]); 
    assign layer_0[2729] = in[91]; 
    assign layer_0[2730] = in[139] & ~in[158]; 
    assign layer_0[2731] = in[35] ^ in[182]; 
    assign layer_0[2732] = in[55] & ~in[152]; 
    assign layer_0[2733] = ~(in[79] ^ in[114]); 
    assign layer_0[2734] = ~in[151] | (in[154] & in[151]); 
    assign layer_0[2735] = in[52] | in[118]; 
    assign layer_0[2736] = ~in[251] | (in[251] & in[203]); 
    assign layer_0[2737] = ~(in[169] ^ in[230]); 
    assign layer_0[2738] = in[241] ^ in[12]; 
    assign layer_0[2739] = in[252] & ~in[101]; 
    assign layer_0[2740] = in[236] ^ in[99]; 
    assign layer_0[2741] = ~(in[152] | in[82]); 
    assign layer_0[2742] = ~(in[104] | in[124]); 
    assign layer_0[2743] = ~(in[79] | in[245]); 
    assign layer_0[2744] = ~(in[39] | in[102]); 
    assign layer_0[2745] = in[135] & ~in[52]; 
    assign layer_0[2746] = in[87] ^ in[134]; 
    assign layer_0[2747] = ~in[115] | (in[199] & in[115]); 
    assign layer_0[2748] = ~(in[22] ^ in[36]); 
    assign layer_0[2749] = in[171]; 
    assign layer_0[2750] = in[179] ^ in[149]; 
    assign layer_0[2751] = ~(in[26] | in[88]); 
    assign layer_0[2752] = ~(in[132] | in[197]); 
    assign layer_0[2753] = in[123] & ~in[90]; 
    assign layer_0[2754] = in[164] ^ in[182]; 
    assign layer_0[2755] = in[109] ^ in[138]; 
    assign layer_0[2756] = ~(in[91] ^ in[89]); 
    assign layer_0[2757] = ~in[218] | (in[166] & in[218]); 
    assign layer_0[2758] = ~(in[207] ^ in[222]); 
    assign layer_0[2759] = ~(in[25] ^ in[72]); 
    assign layer_0[2760] = in[72] | in[41]; 
    assign layer_0[2761] = in[53] & ~in[9]; 
    assign layer_0[2762] = in[121] | in[5]; 
    assign layer_0[2763] = in[103] ^ in[73]; 
    assign layer_0[2764] = in[22] | in[136]; 
    assign layer_0[2765] = in[45] | in[8]; 
    assign layer_0[2766] = ~in[139]; 
    assign layer_0[2767] = ~(in[177] | in[169]); 
    assign layer_0[2768] = ~(in[205] | in[175]); 
    assign layer_0[2769] = ~in[253]; 
    assign layer_0[2770] = ~in[193] | (in[193] & in[148]); 
    assign layer_0[2771] = ~(in[175] ^ in[143]); 
    assign layer_0[2772] = in[142] | in[62]; 
    assign layer_0[2773] = ~(in[172] | in[74]); 
    assign layer_0[2774] = ~(in[105] ^ in[152]); 
    assign layer_0[2775] = in[115]; 
    assign layer_0[2776] = in[86] | in[54]; 
    assign layer_0[2777] = in[83] ^ in[202]; 
    assign layer_0[2778] = ~in[151] | (in[68] & in[151]); 
    assign layer_0[2779] = ~(in[178] ^ in[180]); 
    assign layer_0[2780] = in[69] ^ in[52]; 
    assign layer_0[2781] = ~(in[205] | in[173]); 
    assign layer_0[2782] = in[99] ^ in[41]; 
    assign layer_0[2783] = ~in[25] | (in[87] & in[25]); 
    assign layer_0[2784] = ~in[135] | (in[135] & in[140]); 
    assign layer_0[2785] = ~(in[39] ^ in[181]); 
    assign layer_0[2786] = ~in[40] | (in[40] & in[149]); 
    assign layer_0[2787] = ~(in[112] | in[156]); 
    assign layer_0[2788] = 1'b1; 
    assign layer_0[2789] = in[217] | in[202]; 
    assign layer_0[2790] = ~(in[150] | in[83]); 
    assign layer_0[2791] = in[182] ^ in[180]; 
    assign layer_0[2792] = in[93] | in[86]; 
    assign layer_0[2793] = ~(in[203] | in[23]); 
    assign layer_0[2794] = in[72] ^ in[107]; 
    assign layer_0[2795] = in[83] ^ in[179]; 
    assign layer_0[2796] = ~(in[185] ^ in[247]); 
    assign layer_0[2797] = in[92] & ~in[59]; 
    assign layer_0[2798] = in[67] | in[155]; 
    assign layer_0[2799] = in[228]; 
    assign layer_0[2800] = ~in[105] | (in[105] & in[202]); 
    assign layer_0[2801] = in[24] & ~in[149]; 
    assign layer_0[2802] = in[72] ^ in[210]; 
    assign layer_0[2803] = in[145] | in[120]; 
    assign layer_0[2804] = in[108]; 
    assign layer_0[2805] = ~(in[182] | in[180]); 
    assign layer_0[2806] = in[243] | in[22]; 
    assign layer_0[2807] = in[172] ^ in[72]; 
    assign layer_0[2808] = in[50] | in[209]; 
    assign layer_0[2809] = in[115] | in[30]; 
    assign layer_0[2810] = in[52] ^ in[98]; 
    assign layer_0[2811] = in[137] ^ in[215]; 
    assign layer_0[2812] = ~(in[29] | in[251]); 
    assign layer_0[2813] = in[106] & ~in[72]; 
    assign layer_0[2814] = in[56] & ~in[244]; 
    assign layer_0[2815] = in[121] ^ in[114]; 
    assign layer_0[2816] = in[44] & ~in[22]; 
    assign layer_0[2817] = in[54] | in[69]; 
    assign layer_0[2818] = in[172]; 
    assign layer_0[2819] = in[74] & ~in[120]; 
    assign layer_0[2820] = ~(in[154] | in[131]); 
    assign layer_0[2821] = ~in[73] | (in[73] & in[126]); 
    assign layer_0[2822] = in[135] & in[140]; 
    assign layer_0[2823] = in[153] & ~in[132]; 
    assign layer_0[2824] = in[58]; 
    assign layer_0[2825] = ~(in[233] | in[216]); 
    assign layer_0[2826] = ~in[157]; 
    assign layer_0[2827] = in[180] ^ in[151]; 
    assign layer_0[2828] = in[77] | in[69]; 
    assign layer_0[2829] = ~(in[147] | in[103]); 
    assign layer_0[2830] = ~in[148]; 
    assign layer_0[2831] = ~(in[87] ^ in[107]); 
    assign layer_0[2832] = ~(in[122] | in[23]); 
    assign layer_0[2833] = in[133] | in[135]; 
    assign layer_0[2834] = in[107] & ~in[201]; 
    assign layer_0[2835] = in[89] ^ in[232]; 
    assign layer_0[2836] = in[229] & ~in[149]; 
    assign layer_0[2837] = ~(in[36] | in[81]); 
    assign layer_0[2838] = ~(in[75] ^ in[93]); 
    assign layer_0[2839] = ~(in[85] | in[164]); 
    assign layer_0[2840] = ~in[154] | (in[154] & in[229]); 
    assign layer_0[2841] = in[134] & ~in[53]; 
    assign layer_0[2842] = ~(in[37] | in[210]); 
    assign layer_0[2843] = in[106] ^ in[125]; 
    assign layer_0[2844] = ~in[91] | (in[91] & in[198]); 
    assign layer_0[2845] = in[107] | in[230]; 
    assign layer_0[2846] = in[87] | in[78]; 
    assign layer_0[2847] = ~(in[166] | in[74]); 
    assign layer_0[2848] = in[19]; 
    assign layer_0[2849] = in[131] | in[129]; 
    assign layer_0[2850] = ~in[75] | (in[138] & in[75]); 
    assign layer_0[2851] = ~(in[206] | in[40]); 
    assign layer_0[2852] = ~in[184] | (in[196] & in[184]); 
    assign layer_0[2853] = in[241] | in[20]; 
    assign layer_0[2854] = in[73] ^ in[28]; 
    assign layer_0[2855] = ~(in[151] ^ in[181]); 
    assign layer_0[2856] = in[165]; 
    assign layer_0[2857] = ~(in[131] ^ in[149]); 
    assign layer_0[2858] = in[186] ^ in[166]; 
    assign layer_0[2859] = ~(in[42] | in[37]); 
    assign layer_0[2860] = ~(in[250] ^ in[247]); 
    assign layer_0[2861] = ~(in[101] ^ in[98]); 
    assign layer_0[2862] = ~(in[108] ^ in[90]); 
    assign layer_0[2863] = in[122]; 
    assign layer_0[2864] = ~in[138] | (in[204] & in[138]); 
    assign layer_0[2865] = in[237] | in[169]; 
    assign layer_0[2866] = in[250] ^ in[236]; 
    assign layer_0[2867] = in[165] & ~in[22]; 
    assign layer_0[2868] = ~(in[182] | in[180]); 
    assign layer_0[2869] = in[52] & ~in[99]; 
    assign layer_0[2870] = ~in[76] | (in[76] & in[117]); 
    assign layer_0[2871] = ~(in[37] ^ in[89]); 
    assign layer_0[2872] = in[217] | in[252]; 
    assign layer_0[2873] = ~(in[147] ^ in[206]); 
    assign layer_0[2874] = ~(in[118] | in[245]); 
    assign layer_0[2875] = ~in[86] | (in[86] & in[171]); 
    assign layer_0[2876] = in[232] ^ in[197]; 
    assign layer_0[2877] = ~(in[180] ^ in[181]); 
    assign layer_0[2878] = ~in[120] | (in[120] & in[188]); 
    assign layer_0[2879] = ~(in[108] ^ in[90]); 
    assign layer_0[2880] = ~(in[178] | in[40]); 
    assign layer_0[2881] = in[53] ^ in[22]; 
    assign layer_0[2882] = in[184] | in[153]; 
    assign layer_0[2883] = ~(in[203] | in[21]); 
    assign layer_0[2884] = ~(in[85] | in[106]); 
    assign layer_0[2885] = ~(in[148] | in[113]); 
    assign layer_0[2886] = ~in[132]; 
    assign layer_0[2887] = ~(in[199] ^ in[36]); 
    assign layer_0[2888] = in[120] & ~in[165]; 
    assign layer_0[2889] = ~(in[148] ^ in[166]); 
    assign layer_0[2890] = ~in[155]; 
    assign layer_0[2891] = in[182] ^ in[200]; 
    assign layer_0[2892] = ~(in[247] ^ in[119]); 
    assign layer_0[2893] = ~in[7] | (in[123] & in[7]); 
    assign layer_0[2894] = ~in[149]; 
    assign layer_0[2895] = in[171] ^ in[173]; 
    assign layer_0[2896] = ~in[119]; 
    assign layer_0[2897] = in[72]; 
    assign layer_0[2898] = ~(in[185] ^ in[232]); 
    assign layer_0[2899] = ~in[68]; 
    assign layer_0[2900] = in[220]; 
    assign layer_0[2901] = ~(in[26] ^ in[184]); 
    assign layer_0[2902] = in[4] | in[193]; 
    assign layer_0[2903] = in[148] & ~in[120]; 
    assign layer_0[2904] = in[75] & ~in[87]; 
    assign layer_0[2905] = in[141] & ~in[61]; 
    assign layer_0[2906] = ~in[171] | (in[171] & in[121]); 
    assign layer_0[2907] = in[183] ^ in[121]; 
    assign layer_0[2908] = in[243] | in[171]; 
    assign layer_0[2909] = in[91] | in[89]; 
    assign layer_0[2910] = in[203] ^ in[234]; 
    assign layer_0[2911] = in[125] ^ in[107]; 
    assign layer_0[2912] = in[23] | in[76]; 
    assign layer_0[2913] = ~(in[183] | in[63]); 
    assign layer_0[2914] = ~(in[115] ^ in[133]); 
    assign layer_0[2915] = in[51] ^ in[47]; 
    assign layer_0[2916] = ~(in[146] | in[200]); 
    assign layer_0[2917] = in[131] | in[129]; 
    assign layer_0[2918] = in[164] ^ in[198]; 
    assign layer_0[2919] = ~(in[141] | in[58]); 
    assign layer_0[2920] = ~(in[83] | in[109]); 
    assign layer_0[2921] = in[203]; 
    assign layer_0[2922] = ~(in[44] | in[248]); 
    assign layer_0[2923] = in[131] | in[20]; 
    assign layer_0[2924] = ~in[138]; 
    assign layer_0[2925] = in[53] ^ in[89]; 
    assign layer_0[2926] = in[71] ^ in[213]; 
    assign layer_0[2927] = ~(in[130] ^ in[117]); 
    assign layer_0[2928] = in[147] & ~in[43]; 
    assign layer_0[2929] = ~(in[245] | in[194]); 
    assign layer_0[2930] = in[106] & ~in[186]; 
    assign layer_0[2931] = ~(in[139] | in[103]); 
    assign layer_0[2932] = in[40] ^ in[56]; 
    assign layer_0[2933] = ~in[54] | (in[54] & in[137]); 
    assign layer_0[2934] = ~(in[103] ^ in[72]); 
    assign layer_0[2935] = ~in[119] | (in[82] & in[119]); 
    assign layer_0[2936] = in[55] & in[103]; 
    assign layer_0[2937] = in[210] & ~in[200]; 
    assign layer_0[2938] = ~(in[213] ^ in[244]); 
    assign layer_0[2939] = in[199] ^ in[45]; 
    assign layer_0[2940] = ~(in[53] ^ in[216]); 
    assign layer_0[2941] = ~in[90] | (in[90] & in[28]); 
    assign layer_0[2942] = ~(in[67] ^ in[36]); 
    assign layer_0[2943] = ~in[141] | (in[141] & in[197]); 
    assign layer_0[2944] = ~(in[87] ^ in[39]); 
    assign layer_0[2945] = in[244] & ~in[216]; 
    assign layer_0[2946] = ~in[137]; 
    assign layer_0[2947] = in[98] | in[59]; 
    assign layer_0[2948] = ~(in[131] | in[148]); 
    assign layer_0[2949] = in[93]; 
    assign layer_0[2950] = ~(in[205] | in[28]); 
    assign layer_0[2951] = in[166] | in[120]; 
    assign layer_0[2952] = ~(in[167] | in[151]); 
    assign layer_0[2953] = ~(in[151] | in[60]); 
    assign layer_0[2954] = ~in[140] | (in[59] & in[140]); 
    assign layer_0[2955] = in[196] ^ in[242]; 
    assign layer_0[2956] = in[213] | in[215]; 
    assign layer_0[2957] = in[87] ^ in[228]; 
    assign layer_0[2958] = in[172] ^ in[174]; 
    assign layer_0[2959] = ~(in[43] ^ in[199]); 
    assign layer_0[2960] = in[246] & ~in[214]; 
    assign layer_0[2961] = in[168] & ~in[39]; 
    assign layer_0[2962] = ~(in[157] ^ in[188]); 
    assign layer_0[2963] = in[92]; 
    assign layer_0[2964] = ~(in[65] ^ in[46]); 
    assign layer_0[2965] = in[44] & in[109]; 
    assign layer_0[2966] = in[79] ^ in[93]; 
    assign layer_0[2967] = ~(in[234] ^ in[198]); 
    assign layer_0[2968] = in[116] ^ in[102]; 
    assign layer_0[2969] = ~in[47]; 
    assign layer_0[2970] = ~(in[47] | in[130]); 
    assign layer_0[2971] = ~(in[124] ^ in[156]); 
    assign layer_0[2972] = in[58] | in[42]; 
    assign layer_0[2973] = in[183] & ~in[249]; 
    assign layer_0[2974] = in[192] | in[225]; 
    assign layer_0[2975] = in[178] ^ in[199]; 
    assign layer_0[2976] = in[26] | in[178]; 
    assign layer_0[2977] = ~in[136] | (in[177] & in[136]); 
    assign layer_0[2978] = in[228] ^ in[197]; 
    assign layer_0[2979] = in[61] ^ in[85]; 
    assign layer_0[2980] = ~(in[180] | in[222]); 
    assign layer_0[2981] = ~in[91]; 
    assign layer_0[2982] = ~in[226] | (in[181] & in[226]); 
    assign layer_0[2983] = in[252] | in[137]; 
    assign layer_0[2984] = in[216] ^ in[249]; 
    assign layer_0[2985] = ~(in[154] ^ in[171]); 
    assign layer_0[2986] = ~(in[243] | in[171]); 
    assign layer_0[2987] = ~(in[248] ^ in[12]); 
    assign layer_0[2988] = ~in[39] | (in[166] & in[39]); 
    assign layer_0[2989] = ~(in[168] ^ in[251]); 
    assign layer_0[2990] = in[100] ^ in[165]; 
    assign layer_0[2991] = ~(in[211] | in[233]); 
    assign layer_0[2992] = in[168]; 
    assign layer_0[2993] = in[207] | in[23]; 
    assign layer_0[2994] = ~in[109]; 
    assign layer_0[2995] = ~(in[168] | in[131]); 
    assign layer_0[2996] = ~(in[95] | in[233]); 
    assign layer_0[2997] = ~(in[183] | in[181]); 
    assign layer_0[2998] = ~in[155] | (in[149] & in[155]); 
    assign layer_0[2999] = in[76] & ~in[122]; 
    assign layer_0[3000] = in[61] | in[162]; 
    assign layer_0[3001] = ~(in[154] & in[138]); 
    assign layer_0[3002] = in[39] | in[212]; 
    assign layer_0[3003] = in[92] ^ in[90]; 
    assign layer_0[3004] = in[155] | in[99]; 
    assign layer_0[3005] = in[70]; 
    assign layer_0[3006] = in[53] | in[67]; 
    assign layer_0[3007] = ~(in[215] ^ in[186]); 
    assign layer_0[3008] = ~in[151] | (in[151] & in[117]); 
    assign layer_0[3009] = in[166]; 
    assign layer_0[3010] = ~(in[21] ^ in[51]); 
    assign layer_0[3011] = in[152] & ~in[100]; 
    assign layer_0[3012] = ~(in[210] ^ in[69]); 
    assign layer_0[3013] = ~(in[151] ^ in[120]); 
    assign layer_0[3014] = in[251] ^ in[138]; 
    assign layer_0[3015] = ~(in[243] | in[149]); 
    assign layer_0[3016] = in[98]; 
    assign layer_0[3017] = ~(in[97] ^ in[130]); 
    assign layer_0[3018] = in[197] | in[179]; 
    assign layer_0[3019] = ~in[230] | (in[230] & in[155]); 
    assign layer_0[3020] = ~in[53] | (in[53] & in[148]); 
    assign layer_0[3021] = in[244]; 
    assign layer_0[3022] = ~(in[164] ^ in[181]); 
    assign layer_0[3023] = in[194] ^ in[135]; 
    assign layer_0[3024] = in[248] ^ in[230]; 
    assign layer_0[3025] = in[40] | in[56]; 
    assign layer_0[3026] = ~(in[29] | in[11]); 
    assign layer_0[3027] = in[120] & ~in[140]; 
    assign layer_0[3028] = ~(in[92] ^ in[88]); 
    assign layer_0[3029] = ~(in[21] ^ in[27]); 
    assign layer_0[3030] = in[44] ^ in[91]; 
    assign layer_0[3031] = ~(in[52] | in[57]); 
    assign layer_0[3032] = in[150] & in[149]; 
    assign layer_0[3033] = ~in[58]; 
    assign layer_0[3034] = ~(in[35] | in[150]); 
    assign layer_0[3035] = ~(in[130] | in[58]); 
    assign layer_0[3036] = in[43] | in[108]; 
    assign layer_0[3037] = ~(in[183] ^ in[88]); 
    assign layer_0[3038] = in[182] ^ in[228]; 
    assign layer_0[3039] = in[184] & ~in[60]; 
    assign layer_0[3040] = in[163] ^ in[67]; 
    assign layer_0[3041] = in[103] & ~in[71]; 
    assign layer_0[3042] = in[205] ^ in[178]; 
    assign layer_0[3043] = ~(in[102] ^ in[56]); 
    assign layer_0[3044] = ~(in[163] | in[183]); 
    assign layer_0[3045] = in[73] & ~in[213]; 
    assign layer_0[3046] = ~(in[107] | in[99]); 
    assign layer_0[3047] = ~(in[139] ^ in[213]); 
    assign layer_0[3048] = in[83] ^ in[101]; 
    assign layer_0[3049] = ~(in[9] | in[27]); 
    assign layer_0[3050] = in[157] | in[140]; 
    assign layer_0[3051] = ~(in[131] | in[171]); 
    assign layer_0[3052] = in[172] | in[131]; 
    assign layer_0[3053] = in[120] | in[34]; 
    assign layer_0[3054] = ~(in[149] | in[40]); 
    assign layer_0[3055] = ~in[101] | (in[101] & in[141]); 
    assign layer_0[3056] = in[162] ^ in[62]; 
    assign layer_0[3057] = ~(in[113] ^ in[123]); 
    assign layer_0[3058] = in[106] ^ in[58]; 
    assign layer_0[3059] = ~(in[201] ^ in[198]); 
    assign layer_0[3060] = in[107] | in[75]; 
    assign layer_0[3061] = ~in[137] | (in[137] & in[171]); 
    assign layer_0[3062] = ~(in[172] ^ in[88]); 
    assign layer_0[3063] = in[55]; 
    assign layer_0[3064] = ~(in[60] ^ in[189]); 
    assign layer_0[3065] = in[210] ^ in[245]; 
    assign layer_0[3066] = in[54] & ~in[102]; 
    assign layer_0[3067] = ~(in[111] | in[109]); 
    assign layer_0[3068] = in[139] | in[120]; 
    assign layer_0[3069] = ~in[73] | (in[195] & in[73]); 
    assign layer_0[3070] = in[237] ^ in[205]; 
    assign layer_0[3071] = in[187] ^ in[232]; 
    assign layer_0[3072] = in[214] ^ in[246]; 
    assign layer_0[3073] = ~(in[154] & in[150]); 
    assign layer_0[3074] = ~(in[180] ^ in[182]); 
    assign layer_0[3075] = ~(in[174] | in[157]); 
    assign layer_0[3076] = in[165] | in[118]; 
    assign layer_0[3077] = ~(in[245] | in[248]); 
    assign layer_0[3078] = ~(in[118] ^ in[132]); 
    assign layer_0[3079] = ~in[213] | (in[213] & in[86]); 
    assign layer_0[3080] = in[20] | in[69]; 
    assign layer_0[3081] = ~(in[78] | in[162]); 
    assign layer_0[3082] = ~(in[106] ^ in[103]); 
    assign layer_0[3083] = ~(in[4] | in[95]); 
    assign layer_0[3084] = ~(in[211] ^ in[219]); 
    assign layer_0[3085] = in[114] ^ in[100]; 
    assign layer_0[3086] = ~(in[52] | in[74]); 
    assign layer_0[3087] = in[126] | in[125]; 
    assign layer_0[3088] = ~in[57] | (in[194] & in[57]); 
    assign layer_0[3089] = in[181]; 
    assign layer_0[3090] = in[105]; 
    assign layer_0[3091] = in[147]; 
    assign layer_0[3092] = ~in[89]; 
    assign layer_0[3093] = in[166] ^ in[244]; 
    assign layer_0[3094] = ~in[210]; 
    assign layer_0[3095] = in[78] ^ in[54]; 
    assign layer_0[3096] = in[161] | in[163]; 
    assign layer_0[3097] = in[164] ^ in[199]; 
    assign layer_0[3098] = in[241] ^ in[89]; 
    assign layer_0[3099] = ~(in[206] | in[130]); 
    assign layer_0[3100] = ~in[101]; 
    assign layer_0[3101] = in[130] ^ in[82]; 
    assign layer_0[3102] = ~in[132] | (in[132] & in[122]); 
    assign layer_0[3103] = ~in[173]; 
    assign layer_0[3104] = in[132] | in[88]; 
    assign layer_0[3105] = in[247]; 
    assign layer_0[3106] = in[114] ^ in[85]; 
    assign layer_0[3107] = ~(in[149] | in[146]); 
    assign layer_0[3108] = in[111] | in[205]; 
    assign layer_0[3109] = in[186] & ~in[233]; 
    assign layer_0[3110] = in[132] ^ in[141]; 
    assign layer_0[3111] = ~(in[119] ^ in[150]); 
    assign layer_0[3112] = ~(in[56] ^ in[109]); 
    assign layer_0[3113] = in[21] ^ in[154]; 
    assign layer_0[3114] = in[214]; 
    assign layer_0[3115] = in[222] ^ in[190]; 
    assign layer_0[3116] = ~(in[246] | in[85]); 
    assign layer_0[3117] = in[44] | in[59]; 
    assign layer_0[3118] = ~in[75] | (in[75] & in[118]); 
    assign layer_0[3119] = ~(in[196] ^ in[187]); 
    assign layer_0[3120] = in[27] & ~in[89]; 
    assign layer_0[3121] = in[199] & ~in[120]; 
    assign layer_0[3122] = ~(in[45] | in[63]); 
    assign layer_0[3123] = in[98] | in[38]; 
    assign layer_0[3124] = in[90] & ~in[26]; 
    assign layer_0[3125] = in[7] ^ in[34]; 
    assign layer_0[3126] = in[164] ^ in[182]; 
    assign layer_0[3127] = in[152] & ~in[40]; 
    assign layer_0[3128] = in[110] ^ in[92]; 
    assign layer_0[3129] = ~(in[163] ^ in[194]); 
    assign layer_0[3130] = in[151] & ~in[113]; 
    assign layer_0[3131] = in[141] | in[230]; 
    assign layer_0[3132] = ~(in[157] | in[161]); 
    assign layer_0[3133] = ~(in[94] | in[24]); 
    assign layer_0[3134] = ~(in[134] | in[215]); 
    assign layer_0[3135] = in[79] ^ in[141]; 
    assign layer_0[3136] = in[152] ^ in[89]; 
    assign layer_0[3137] = ~in[236]; 
    assign layer_0[3138] = ~(in[129] ^ in[115]); 
    assign layer_0[3139] = ~(in[119] | in[102]); 
    assign layer_0[3140] = ~(in[104] ^ in[78]); 
    assign layer_0[3141] = in[71] | in[103]; 
    assign layer_0[3142] = in[231] ^ in[171]; 
    assign layer_0[3143] = in[118] ^ in[169]; 
    assign layer_0[3144] = ~in[220] | (in[220] & in[76]); 
    assign layer_0[3145] = in[40] ^ in[75]; 
    assign layer_0[3146] = ~(in[245] ^ in[137]); 
    assign layer_0[3147] = ~in[101]; 
    assign layer_0[3148] = in[197] | in[195]; 
    assign layer_0[3149] = ~(in[8] | in[11]); 
    assign layer_0[3150] = ~(in[121] ^ in[186]); 
    assign layer_0[3151] = in[57] & ~in[180]; 
    assign layer_0[3152] = ~in[57]; 
    assign layer_0[3153] = ~in[138] | (in[138] & in[178]); 
    assign layer_0[3154] = ~(in[97] | in[234]); 
    assign layer_0[3155] = ~(in[103] ^ in[194]); 
    assign layer_0[3156] = ~in[153]; 
    assign layer_0[3157] = in[55]; 
    assign layer_0[3158] = in[78] | in[237]; 
    assign layer_0[3159] = in[88] ^ in[57]; 
    assign layer_0[3160] = in[35] ^ in[125]; 
    assign layer_0[3161] = ~(in[187] ^ in[204]); 
    assign layer_0[3162] = ~in[155] | (in[196] & in[155]); 
    assign layer_0[3163] = in[227] | in[212]; 
    assign layer_0[3164] = in[83] | in[190]; 
    assign layer_0[3165] = in[93] ^ in[70]; 
    assign layer_0[3166] = ~(in[165] ^ in[147]); 
    assign layer_0[3167] = ~(in[63] ^ in[234]); 
    assign layer_0[3168] = ~in[163]; 
    assign layer_0[3169] = in[108] ^ in[90]; 
    assign layer_0[3170] = ~(in[89] ^ in[58]); 
    assign layer_0[3171] = in[63] ^ in[11]; 
    assign layer_0[3172] = in[54] & ~in[116]; 
    assign layer_0[3173] = in[140] | in[122]; 
    assign layer_0[3174] = ~(in[30] | in[79]); 
    assign layer_0[3175] = ~in[212] | (in[231] & in[212]); 
    assign layer_0[3176] = ~(in[218] | in[233]); 
    assign layer_0[3177] = ~in[170] | (in[221] & in[170]); 
    assign layer_0[3178] = ~(in[23] ^ in[58]); 
    assign layer_0[3179] = ~in[206]; 
    assign layer_0[3180] = ~in[9] | (in[43] & in[9]); 
    assign layer_0[3181] = ~(in[213] ^ in[150]); 
    assign layer_0[3182] = ~(in[73] & in[202]); 
    assign layer_0[3183] = in[250] ^ in[165]; 
    assign layer_0[3184] = ~in[228] | (in[228] & in[158]); 
    assign layer_0[3185] = in[204] | in[180]; 
    assign layer_0[3186] = in[47]; 
    assign layer_0[3187] = ~(in[151] & in[121]); 
    assign layer_0[3188] = ~in[76] | (in[76] & in[151]); 
    assign layer_0[3189] = in[199] & ~in[245]; 
    assign layer_0[3190] = ~(in[59] ^ in[88]); 
    assign layer_0[3191] = in[30] ^ in[79]; 
    assign layer_0[3192] = in[163] ^ in[211]; 
    assign layer_0[3193] = in[136] & ~in[141]; 
    assign layer_0[3194] = ~in[222]; 
    assign layer_0[3195] = in[177] ^ in[111]; 
    assign layer_0[3196] = in[131] & ~in[150]; 
    assign layer_0[3197] = ~in[108] | (in[218] & in[108]); 
    assign layer_0[3198] = in[36] ^ in[86]; 
    assign layer_0[3199] = ~(in[163] ^ in[167]); 
    assign layer_0[3200] = in[249] ^ in[233]; 
    assign layer_0[3201] = ~(in[202] ^ in[36]); 
    assign layer_0[3202] = in[139] ^ in[183]; 
    assign layer_0[3203] = ~in[131]; 
    assign layer_0[3204] = in[216] | in[248]; 
    assign layer_0[3205] = in[197] ^ in[169]; 
    assign layer_0[3206] = in[30]; 
    assign layer_0[3207] = in[242] ^ in[141]; 
    assign layer_0[3208] = ~(in[189] ^ in[115]); 
    assign layer_0[3209] = in[122] | in[249]; 
    assign layer_0[3210] = ~(in[150] | in[142]); 
    assign layer_0[3211] = ~(in[136] ^ in[164]); 
    assign layer_0[3212] = in[8] ^ in[10]; 
    assign layer_0[3213] = in[29] ^ in[126]; 
    assign layer_0[3214] = ~in[39]; 
    assign layer_0[3215] = ~in[105]; 
    assign layer_0[3216] = in[109] ^ in[102]; 
    assign layer_0[3217] = in[247] ^ in[249]; 
    assign layer_0[3218] = in[167] ^ in[135]; 
    assign layer_0[3219] = in[230] & ~in[21]; 
    assign layer_0[3220] = ~(in[198] | in[158]); 
    assign layer_0[3221] = in[42] | in[242]; 
    assign layer_0[3222] = ~(in[195] ^ in[112]); 
    assign layer_0[3223] = in[132] | in[110]; 
    assign layer_0[3224] = ~(in[175] | in[206]); 
    assign layer_0[3225] = in[165] & ~in[95]; 
    assign layer_0[3226] = in[74] ^ in[77]; 
    assign layer_0[3227] = ~(in[88] | in[210]); 
    assign layer_0[3228] = in[135] & ~in[190]; 
    assign layer_0[3229] = ~(in[98] | in[100]); 
    assign layer_0[3230] = ~(in[168] | in[166]); 
    assign layer_0[3231] = in[29] ^ in[11]; 
    assign layer_0[3232] = in[92] | in[114]; 
    assign layer_0[3233] = ~(in[181] ^ in[163]); 
    assign layer_0[3234] = in[91] ^ in[73]; 
    assign layer_0[3235] = in[78] | in[199]; 
    assign layer_0[3236] = in[214] | in[245]; 
    assign layer_0[3237] = in[122] & ~in[60]; 
    assign layer_0[3238] = ~in[202] | (in[115] & in[202]); 
    assign layer_0[3239] = in[93] ^ in[91]; 
    assign layer_0[3240] = in[142] | in[245]; 
    assign layer_0[3241] = ~(in[87] ^ in[151]); 
    assign layer_0[3242] = ~(in[184] | in[211]); 
    assign layer_0[3243] = in[132] ^ in[134]; 
    assign layer_0[3244] = in[123] ^ in[154]; 
    assign layer_0[3245] = in[142]; 
    assign layer_0[3246] = in[43] ^ in[79]; 
    assign layer_0[3247] = in[95] ^ in[106]; 
    assign layer_0[3248] = ~(in[74] ^ in[94]); 
    assign layer_0[3249] = ~(in[172] | in[180]); 
    assign layer_0[3250] = ~in[230] | (in[92] & in[230]); 
    assign layer_0[3251] = ~in[221]; 
    assign layer_0[3252] = ~(in[205] ^ in[150]); 
    assign layer_0[3253] = in[231] | in[247]; 
    assign layer_0[3254] = ~(in[106] ^ in[108]); 
    assign layer_0[3255] = ~(in[245] | in[65]); 
    assign layer_0[3256] = ~in[88] | (in[88] & in[84]); 
    assign layer_0[3257] = ~(in[73] ^ in[41]); 
    assign layer_0[3258] = ~(in[230] | in[246]); 
    assign layer_0[3259] = in[145] | in[159]; 
    assign layer_0[3260] = in[100] ^ in[183]; 
    assign layer_0[3261] = ~in[98]; 
    assign layer_0[3262] = in[52] | in[107]; 
    assign layer_0[3263] = in[105] ^ in[72]; 
    assign layer_0[3264] = in[31] | in[20]; 
    assign layer_0[3265] = ~(in[90] ^ in[59]); 
    assign layer_0[3266] = ~(in[92] ^ in[131]); 
    assign layer_0[3267] = ~in[132] | (in[132] & in[206]); 
    assign layer_0[3268] = in[138] | in[72]; 
    assign layer_0[3269] = ~(in[137] ^ in[139]); 
    assign layer_0[3270] = ~in[211]; 
    assign layer_0[3271] = in[85] ^ in[99]; 
    assign layer_0[3272] = in[134] ^ in[143]; 
    assign layer_0[3273] = in[234] ^ in[60]; 
    assign layer_0[3274] = ~(in[119] | in[234]); 
    assign layer_0[3275] = ~(in[195] | in[215]); 
    assign layer_0[3276] = in[70] & ~in[227]; 
    assign layer_0[3277] = in[241] | in[101]; 
    assign layer_0[3278] = ~(in[159] ^ in[211]); 
    assign layer_0[3279] = in[70] ^ in[38]; 
    assign layer_0[3280] = ~(in[116] | in[22]); 
    assign layer_0[3281] = ~(in[132] | in[84]); 
    assign layer_0[3282] = in[181]; 
    assign layer_0[3283] = in[204] & ~in[216]; 
    assign layer_0[3284] = ~in[140] | (in[140] & in[154]); 
    assign layer_0[3285] = in[164] | in[103]; 
    assign layer_0[3286] = in[67] | in[84]; 
    assign layer_0[3287] = in[15] | in[92]; 
    assign layer_0[3288] = in[40] | in[247]; 
    assign layer_0[3289] = in[38] | in[69]; 
    assign layer_0[3290] = in[150] | in[41]; 
    assign layer_0[3291] = in[95] | in[234]; 
    assign layer_0[3292] = in[143]; 
    assign layer_0[3293] = in[58] & ~in[237]; 
    assign layer_0[3294] = ~(in[175] ^ in[206]); 
    assign layer_0[3295] = in[245] & ~in[141]; 
    assign layer_0[3296] = ~(in[149] | in[244]); 
    assign layer_0[3297] = ~in[110]; 
    assign layer_0[3298] = in[148] ^ in[146]; 
    assign layer_0[3299] = in[196] ^ in[178]; 
    assign layer_0[3300] = ~in[202] | (in[202] & in[182]); 
    assign layer_0[3301] = in[167] & ~in[93]; 
    assign layer_0[3302] = ~in[109]; 
    assign layer_0[3303] = in[236] | in[235]; 
    assign layer_0[3304] = ~(in[34] ^ in[117]); 
    assign layer_0[3305] = ~(in[104] ^ in[123]); 
    assign layer_0[3306] = in[184] & ~in[247]; 
    assign layer_0[3307] = in[118] ^ in[104]; 
    assign layer_0[3308] = in[59]; 
    assign layer_0[3309] = ~(in[206] ^ in[136]); 
    assign layer_0[3310] = in[137] ^ in[162]; 
    assign layer_0[3311] = in[59] & ~in[103]; 
    assign layer_0[3312] = ~(in[171] ^ in[156]); 
    assign layer_0[3313] = ~(in[135] ^ in[104]); 
    assign layer_0[3314] = ~(in[99] ^ in[102]); 
    assign layer_0[3315] = ~in[134] | (in[204] & in[134]); 
    assign layer_0[3316] = ~in[242] | (in[203] & in[242]); 
    assign layer_0[3317] = in[186] | in[155]; 
    assign layer_0[3318] = in[235] | in[199]; 
    assign layer_0[3319] = in[94]; 
    assign layer_0[3320] = ~(in[99] & in[83]); 
    assign layer_0[3321] = in[148] ^ in[39]; 
    assign layer_0[3322] = ~in[119] | (in[119] & in[131]); 
    assign layer_0[3323] = in[153]; 
    assign layer_0[3324] = in[231] | in[231]; 
    assign layer_0[3325] = ~(in[217] ^ in[250]); 
    assign layer_0[3326] = in[72] & ~in[138]; 
    assign layer_0[3327] = in[138]; 
    assign layer_0[3328] = in[166] | in[147]; 
    assign layer_0[3329] = ~(in[229] ^ in[56]); 
    assign layer_0[3330] = in[186] & ~in[152]; 
    assign layer_0[3331] = ~(in[231] ^ in[54]); 
    assign layer_0[3332] = ~in[231] | (in[168] & in[231]); 
    assign layer_0[3333] = ~(in[103] ^ in[170]); 
    assign layer_0[3334] = in[73] & ~in[111]; 
    assign layer_0[3335] = ~(in[99] | in[71]); 
    assign layer_0[3336] = in[75] ^ in[116]; 
    assign layer_0[3337] = ~(in[204] | in[106]); 
    assign layer_0[3338] = in[115] ^ in[101]; 
    assign layer_0[3339] = ~(in[90] ^ in[92]); 
    assign layer_0[3340] = ~(in[92] | in[26]); 
    assign layer_0[3341] = in[107] & ~in[74]; 
    assign layer_0[3342] = ~in[236] | (in[236] & in[214]); 
    assign layer_0[3343] = ~(in[77] ^ in[43]); 
    assign layer_0[3344] = ~(in[22] ^ in[70]); 
    assign layer_0[3345] = in[154]; 
    assign layer_0[3346] = ~(in[167] | in[118]); 
    assign layer_0[3347] = ~(in[104] ^ in[212]); 
    assign layer_0[3348] = in[243] ^ in[234]; 
    assign layer_0[3349] = ~(in[152] | in[24]); 
    assign layer_0[3350] = in[214] & ~in[179]; 
    assign layer_0[3351] = in[136] & in[137]; 
    assign layer_0[3352] = in[213] ^ in[211]; 
    assign layer_0[3353] = ~(in[59] ^ in[107]); 
    assign layer_0[3354] = ~(in[52] ^ in[188]); 
    assign layer_0[3355] = ~(in[27] | in[44]); 
    assign layer_0[3356] = in[43] ^ in[53]; 
    assign layer_0[3357] = in[131]; 
    assign layer_0[3358] = in[27] ^ in[106]; 
    assign layer_0[3359] = in[142] ^ in[156]; 
    assign layer_0[3360] = in[105]; 
    assign layer_0[3361] = in[197] | in[235]; 
    assign layer_0[3362] = in[121] & ~in[197]; 
    assign layer_0[3363] = ~(in[41] ^ in[117]); 
    assign layer_0[3364] = ~(in[108] ^ in[110]); 
    assign layer_0[3365] = ~(in[84] ^ in[70]); 
    assign layer_0[3366] = ~(in[139] & in[137]); 
    assign layer_0[3367] = ~in[198] | (in[198] & in[185]); 
    assign layer_0[3368] = ~(in[98] ^ in[167]); 
    assign layer_0[3369] = ~in[130]; 
    assign layer_0[3370] = in[140] ^ in[117]; 
    assign layer_0[3371] = ~(in[176] | in[136]); 
    assign layer_0[3372] = ~(in[105] ^ in[54]); 
    assign layer_0[3373] = ~(in[246] ^ in[215]); 
    assign layer_0[3374] = ~(in[242] | in[251]); 
    assign layer_0[3375] = ~(in[54] ^ in[60]); 
    assign layer_0[3376] = ~in[152] | (in[93] & in[152]); 
    assign layer_0[3377] = ~(in[216] ^ in[187]); 
    assign layer_0[3378] = ~in[165] | (in[165] & in[86]); 
    assign layer_0[3379] = in[213] | in[159]; 
    assign layer_0[3380] = ~in[157]; 
    assign layer_0[3381] = ~in[59]; 
    assign layer_0[3382] = in[99] ^ in[98]; 
    assign layer_0[3383] = in[118]; 
    assign layer_0[3384] = ~in[70]; 
    assign layer_0[3385] = in[163] ^ in[7]; 
    assign layer_0[3386] = ~(in[241] | in[147]); 
    assign layer_0[3387] = in[190] ^ in[86]; 
    assign layer_0[3388] = in[24] ^ in[56]; 
    assign layer_0[3389] = in[152] ^ in[105]; 
    assign layer_0[3390] = in[40]; 
    assign layer_0[3391] = in[51] ^ in[99]; 
    assign layer_0[3392] = in[85] ^ in[155]; 
    assign layer_0[3393] = ~(in[102] ^ in[170]); 
    assign layer_0[3394] = ~in[163] | (in[163] & in[13]); 
    assign layer_0[3395] = in[142] ^ in[46]; 
    assign layer_0[3396] = in[21]; 
    assign layer_0[3397] = in[118] ^ in[88]; 
    assign layer_0[3398] = ~in[97]; 
    assign layer_0[3399] = in[121] | in[170]; 
    assign layer_0[3400] = in[245] & ~in[216]; 
    assign layer_0[3401] = ~(in[205] ^ in[198]); 
    assign layer_0[3402] = ~(in[87] | in[246]); 
    assign layer_0[3403] = in[39] ^ in[87]; 
    assign layer_0[3404] = ~in[200] | (in[42] & in[200]); 
    assign layer_0[3405] = ~in[57] | (in[22] & in[57]); 
    assign layer_0[3406] = in[210] ^ in[245]; 
    assign layer_0[3407] = ~(in[189] ^ in[220]); 
    assign layer_0[3408] = in[113] | in[163]; 
    assign layer_0[3409] = in[135] | in[188]; 
    assign layer_0[3410] = in[102] ^ in[236]; 
    assign layer_0[3411] = in[214] | in[228]; 
    assign layer_0[3412] = in[200] ^ in[52]; 
    assign layer_0[3413] = in[117] ^ in[155]; 
    assign layer_0[3414] = ~in[168] | (in[168] & in[126]); 
    assign layer_0[3415] = in[179] & ~in[160]; 
    assign layer_0[3416] = ~in[54]; 
    assign layer_0[3417] = in[25] | in[190]; 
    assign layer_0[3418] = ~in[167] | (in[167] & in[163]); 
    assign layer_0[3419] = ~(in[31] | in[12]); 
    assign layer_0[3420] = ~(in[241] | in[174]); 
    assign layer_0[3421] = in[88] ^ in[103]; 
    assign layer_0[3422] = in[37] | in[197]; 
    assign layer_0[3423] = ~(in[68] ^ in[204]); 
    assign layer_0[3424] = ~(in[140] | in[75]); 
    assign layer_0[3425] = ~in[152] | (in[152] & in[69]); 
    assign layer_0[3426] = ~(in[55] | in[56]); 
    assign layer_0[3427] = ~(in[173] ^ in[117]); 
    assign layer_0[3428] = in[221] ^ in[190]; 
    assign layer_0[3429] = in[139] | in[113]; 
    assign layer_0[3430] = in[233] | in[146]; 
    assign layer_0[3431] = ~(in[195] ^ in[137]); 
    assign layer_0[3432] = ~in[84]; 
    assign layer_0[3433] = ~(in[42] | in[53]); 
    assign layer_0[3434] = in[25] & in[148]; 
    assign layer_0[3435] = in[141] ^ in[127]; 
    assign layer_0[3436] = ~(in[147] ^ in[133]); 
    assign layer_0[3437] = ~(in[90] ^ in[92]); 
    assign layer_0[3438] = in[209] ^ in[152]; 
    assign layer_0[3439] = ~(in[249] ^ in[219]); 
    assign layer_0[3440] = in[203] | in[202]; 
    assign layer_0[3441] = in[207] | in[9]; 
    assign layer_0[3442] = in[199] ^ in[54]; 
    assign layer_0[3443] = in[101] & ~in[190]; 
    assign layer_0[3444] = ~(in[28] ^ in[47]); 
    assign layer_0[3445] = in[207]; 
    assign layer_0[3446] = in[110] | in[142]; 
    assign layer_0[3447] = ~(in[76] ^ in[44]); 
    assign layer_0[3448] = in[188] | in[21]; 
    assign layer_0[3449] = ~in[136] | (in[5] & in[136]); 
    assign layer_0[3450] = ~(in[150] ^ in[182]); 
    assign layer_0[3451] = in[87] & ~in[212]; 
    assign layer_0[3452] = ~(in[146] | in[118]); 
    assign layer_0[3453] = in[146] | in[164]; 
    assign layer_0[3454] = in[192] | in[11]; 
    assign layer_0[3455] = ~in[75]; 
    assign layer_0[3456] = ~(in[103] ^ in[134]); 
    assign layer_0[3457] = ~in[121] | (in[121] & in[196]); 
    assign layer_0[3458] = in[28] ^ in[62]; 
    assign layer_0[3459] = ~(in[157] | in[90]); 
    assign layer_0[3460] = ~(in[136] ^ in[181]); 
    assign layer_0[3461] = ~(in[139] ^ in[24]); 
    assign layer_0[3462] = in[107] & ~in[89]; 
    assign layer_0[3463] = in[213] ^ in[211]; 
    assign layer_0[3464] = in[186] & in[221]; 
    assign layer_0[3465] = ~in[87] | (in[87] & in[242]); 
    assign layer_0[3466] = ~in[34]; 
    assign layer_0[3467] = in[57] & ~in[131]; 
    assign layer_0[3468] = in[143] ^ in[190]; 
    assign layer_0[3469] = in[52] & ~in[38]; 
    assign layer_0[3470] = ~(in[66] ^ in[188]); 
    assign layer_0[3471] = ~in[153] | (in[236] & in[153]); 
    assign layer_0[3472] = ~(in[76] | in[91]); 
    assign layer_0[3473] = ~(in[54] | in[38]); 
    assign layer_0[3474] = in[107] & ~in[41]; 
    assign layer_0[3475] = in[88] | in[89]; 
    assign layer_0[3476] = ~(in[40] ^ in[87]); 
    assign layer_0[3477] = in[118] ^ in[133]; 
    assign layer_0[3478] = in[200] ^ in[181]; 
    assign layer_0[3479] = ~in[151]; 
    assign layer_0[3480] = ~(in[103] ^ in[86]); 
    assign layer_0[3481] = in[50] ^ in[82]; 
    assign layer_0[3482] = ~(in[198] ^ in[229]); 
    assign layer_0[3483] = in[63] ^ in[93]; 
    assign layer_0[3484] = in[40] ^ in[72]; 
    assign layer_0[3485] = in[43] | in[58]; 
    assign layer_0[3486] = in[164] | in[90]; 
    assign layer_0[3487] = ~(in[150] ^ in[54]); 
    assign layer_0[3488] = ~(in[130] ^ in[132]); 
    assign layer_0[3489] = in[87] ^ in[39]; 
    assign layer_0[3490] = in[203] ^ in[234]; 
    assign layer_0[3491] = ~in[171] | (in[120] & in[171]); 
    assign layer_0[3492] = in[188] ^ in[250]; 
    assign layer_0[3493] = ~in[8] | (in[42] & in[8]); 
    assign layer_0[3494] = ~(in[75] ^ in[107]); 
    assign layer_0[3495] = in[119] & ~in[187]; 
    assign layer_0[3496] = ~in[161]; 
    assign layer_0[3497] = in[221]; 
    assign layer_0[3498] = in[87] ^ in[88]; 
    assign layer_0[3499] = ~(in[250] ^ in[58]); 
    assign layer_0[3500] = ~in[11]; 
    assign layer_0[3501] = ~(in[111] ^ in[93]); 
    assign layer_0[3502] = ~(in[218] ^ in[187]); 
    assign layer_0[3503] = ~(in[183] ^ in[180]); 
    assign layer_0[3504] = ~(in[12] | in[203]); 
    assign layer_0[3505] = in[124] | in[157]; 
    assign layer_0[3506] = ~(in[52] ^ in[150]); 
    assign layer_0[3507] = in[166] ^ in[132]; 
    assign layer_0[3508] = in[54] ^ in[22]; 
    assign layer_0[3509] = in[88] ^ in[120]; 
    assign layer_0[3510] = ~(in[102] | in[200]); 
    assign layer_0[3511] = in[76] | in[83]; 
    assign layer_0[3512] = in[100] ^ in[86]; 
    assign layer_0[3513] = in[150] ^ in[148]; 
    assign layer_0[3514] = ~(in[165] | in[162]); 
    assign layer_0[3515] = in[73] ^ in[75]; 
    assign layer_0[3516] = ~(in[152] | in[121]); 
    assign layer_0[3517] = in[147] | in[85]; 
    assign layer_0[3518] = ~(in[161] ^ in[169]); 
    assign layer_0[3519] = ~(in[200] ^ in[233]); 
    assign layer_0[3520] = in[230] ^ in[57]; 
    assign layer_0[3521] = ~(in[236] & in[67]); 
    assign layer_0[3522] = in[175] ^ in[243]; 
    assign layer_0[3523] = in[99] ^ in[54]; 
    assign layer_0[3524] = ~(in[117] | in[79]); 
    assign layer_0[3525] = ~(in[113] | in[223]); 
    assign layer_0[3526] = ~(in[215] ^ in[55]); 
    assign layer_0[3527] = ~(in[149] ^ in[147]); 
    assign layer_0[3528] = ~(in[92] ^ in[94]); 
    assign layer_0[3529] = in[107] ^ in[140]; 
    assign layer_0[3530] = in[246] | in[78]; 
    assign layer_0[3531] = ~(in[124] ^ in[231]); 
    assign layer_0[3532] = ~(in[232] ^ in[21]); 
    assign layer_0[3533] = in[76] ^ in[139]; 
    assign layer_0[3534] = in[250]; 
    assign layer_0[3535] = in[92] ^ in[95]; 
    assign layer_0[3536] = in[199] | in[180]; 
    assign layer_0[3537] = in[166]; 
    assign layer_0[3538] = in[70] ^ in[84]; 
    assign layer_0[3539] = ~(in[242] | in[120]); 
    assign layer_0[3540] = in[103] ^ in[117]; 
    assign layer_0[3541] = in[127] ^ in[8]; 
    assign layer_0[3542] = in[251] | in[235]; 
    assign layer_0[3543] = ~(in[132] ^ in[130]); 
    assign layer_0[3544] = ~in[169]; 
    assign layer_0[3545] = ~(in[12] ^ in[9]); 
    assign layer_0[3546] = in[228] ^ in[24]; 
    assign layer_0[3547] = ~in[105]; 
    assign layer_0[3548] = in[50] | in[171]; 
    assign layer_0[3549] = in[82] | in[98]; 
    assign layer_0[3550] = ~(in[132] ^ in[134]); 
    assign layer_0[3551] = ~(in[198] ^ in[61]); 
    assign layer_0[3552] = ~in[95]; 
    assign layer_0[3553] = in[20] & in[56]; 
    assign layer_0[3554] = in[89]; 
    assign layer_0[3555] = ~(in[77] ^ in[75]); 
    assign layer_0[3556] = in[39] & in[174]; 
    assign layer_0[3557] = ~(in[91] ^ in[119]); 
    assign layer_0[3558] = in[121] & ~in[118]; 
    assign layer_0[3559] = ~(in[150] | in[132]); 
    assign layer_0[3560] = in[72] | in[41]; 
    assign layer_0[3561] = ~in[215] | (in[215] & in[150]); 
    assign layer_0[3562] = in[156] ^ in[138]; 
    assign layer_0[3563] = ~(in[55] & in[54]); 
    assign layer_0[3564] = in[156] ^ in[137]; 
    assign layer_0[3565] = in[45] ^ in[79]; 
    assign layer_0[3566] = in[119] & ~in[115]; 
    assign layer_0[3567] = in[36] ^ in[50]; 
    assign layer_0[3568] = ~(in[98] | in[147]); 
    assign layer_0[3569] = ~in[230] | (in[170] & in[230]); 
    assign layer_0[3570] = ~in[169] | (in[20] & in[169]); 
    assign layer_0[3571] = ~(in[53] | in[211]); 
    assign layer_0[3572] = in[12] | in[200]; 
    assign layer_0[3573] = in[138] & ~in[39]; 
    assign layer_0[3574] = ~(in[43] & in[39]); 
    assign layer_0[3575] = in[95] ^ in[61]; 
    assign layer_0[3576] = ~in[199]; 
    assign layer_0[3577] = in[102] ^ in[162]; 
    assign layer_0[3578] = ~(in[237] ^ in[206]); 
    assign layer_0[3579] = ~(in[198] ^ in[146]); 
    assign layer_0[3580] = ~(in[121] ^ in[162]); 
    assign layer_0[3581] = ~in[138]; 
    assign layer_0[3582] = in[86] ^ in[38]; 
    assign layer_0[3583] = in[219] | in[194]; 
    assign layer_0[3584] = in[35] ^ in[66]; 
    assign layer_0[3585] = in[138] ^ in[156]; 
    assign layer_0[3586] = ~(in[165] ^ in[24]); 
    assign layer_0[3587] = in[152] & ~in[108]; 
    assign layer_0[3588] = ~(in[184] & in[72]); 
    assign layer_0[3589] = in[59] ^ in[87]; 
    assign layer_0[3590] = ~(in[125] | in[191]); 
    assign layer_0[3591] = in[198] ^ in[244]; 
    assign layer_0[3592] = ~in[120] | (in[62] & in[120]); 
    assign layer_0[3593] = ~(in[98] | in[99]); 
    assign layer_0[3594] = ~in[216] | (in[216] & in[124]); 
    assign layer_0[3595] = ~(in[147] | in[182]); 
    assign layer_0[3596] = ~(in[70] | in[90]); 
    assign layer_0[3597] = ~in[199] | (in[199] & in[42]); 
    assign layer_0[3598] = ~(in[159] ^ in[141]); 
    assign layer_0[3599] = ~in[149]; 
    assign layer_0[3600] = ~(in[71] | in[245]); 
    assign layer_0[3601] = in[187] & ~in[38]; 
    assign layer_0[3602] = in[249] ^ in[248]; 
    assign layer_0[3603] = ~(in[164] | in[182]); 
    assign layer_0[3604] = in[162] ^ in[249]; 
    assign layer_0[3605] = ~(in[164] ^ in[167]); 
    assign layer_0[3606] = in[116] | in[213]; 
    assign layer_0[3607] = ~in[219] | (in[99] & in[219]); 
    assign layer_0[3608] = in[203] & ~in[81]; 
    assign layer_0[3609] = in[249] ^ in[246]; 
    assign layer_0[3610] = ~(in[118] & in[198]); 
    assign layer_0[3611] = in[142] | in[157]; 
    assign layer_0[3612] = ~in[198] | (in[198] & in[244]); 
    assign layer_0[3613] = ~(in[211] | in[237]); 
    assign layer_0[3614] = in[149]; 
    assign layer_0[3615] = in[244]; 
    assign layer_0[3616] = ~in[153] | (in[203] & in[153]); 
    assign layer_0[3617] = in[141]; 
    assign layer_0[3618] = in[170]; 
    assign layer_0[3619] = ~(in[100] ^ in[114]); 
    assign layer_0[3620] = in[55] ^ in[25]; 
    assign layer_0[3621] = in[81] | in[50]; 
    assign layer_0[3622] = ~(in[168] ^ in[183]); 
    assign layer_0[3623] = ~(in[150] ^ in[76]); 
    assign layer_0[3624] = in[133] | in[142]; 
    assign layer_0[3625] = in[94] ^ in[95]; 
    assign layer_0[3626] = in[202] & ~in[90]; 
    assign layer_0[3627] = ~(in[172] ^ in[242]); 
    assign layer_0[3628] = in[91] ^ in[93]; 
    assign layer_0[3629] = in[120] ^ in[116]; 
    assign layer_0[3630] = ~in[70] | (in[70] & in[26]); 
    assign layer_0[3631] = ~(in[91] | in[92]); 
    assign layer_0[3632] = ~in[197]; 
    assign layer_0[3633] = ~(in[71] | in[57]); 
    assign layer_0[3634] = in[62] | in[196]; 
    assign layer_0[3635] = in[120] ^ in[189]; 
    assign layer_0[3636] = ~(in[123] ^ in[90]); 
    assign layer_0[3637] = in[194] ^ in[213]; 
    assign layer_0[3638] = ~(in[122] ^ in[8]); 
    assign layer_0[3639] = in[44] ^ in[42]; 
    assign layer_0[3640] = ~(in[154] ^ in[20]); 
    assign layer_0[3641] = in[55] ^ in[103]; 
    assign layer_0[3642] = in[53] | in[74]; 
    assign layer_0[3643] = in[173] | in[132]; 
    assign layer_0[3644] = ~(in[250] ^ in[75]); 
    assign layer_0[3645] = in[198] ^ in[229]; 
    assign layer_0[3646] = ~in[152]; 
    assign layer_0[3647] = in[170] ^ in[179]; 
    assign layer_0[3648] = ~(in[92] ^ in[61]); 
    assign layer_0[3649] = in[115] ^ in[117]; 
    assign layer_0[3650] = in[168] & ~in[66]; 
    assign layer_0[3651] = in[197]; 
    assign layer_0[3652] = in[121] ^ in[168]; 
    assign layer_0[3653] = ~(in[149] ^ in[134]); 
    assign layer_0[3654] = in[119] ^ in[69]; 
    assign layer_0[3655] = in[170] ^ in[105]; 
    assign layer_0[3656] = ~(in[148] | in[146]); 
    assign layer_0[3657] = in[20] & ~in[45]; 
    assign layer_0[3658] = ~(in[212] ^ in[249]); 
    assign layer_0[3659] = in[114] ^ in[101]; 
    assign layer_0[3660] = in[221] | in[211]; 
    assign layer_0[3661] = ~(in[221] | in[235]); 
    assign layer_0[3662] = in[5] ^ in[53]; 
    assign layer_0[3663] = in[89] & ~in[8]; 
    assign layer_0[3664] = in[105] | in[34]; 
    assign layer_0[3665] = in[106] & ~in[233]; 
    assign layer_0[3666] = in[217] ^ in[151]; 
    assign layer_0[3667] = ~(in[91] | in[137]); 
    assign layer_0[3668] = in[125] | in[169]; 
    assign layer_0[3669] = in[139] | in[92]; 
    assign layer_0[3670] = ~in[148]; 
    assign layer_0[3671] = in[136] ^ in[22]; 
    assign layer_0[3672] = ~in[71] | (in[130] & in[71]); 
    assign layer_0[3673] = ~in[123] | (in[123] & in[164]); 
    assign layer_0[3674] = in[113] | in[244]; 
    assign layer_0[3675] = ~in[244]; 
    assign layer_0[3676] = ~(in[92] ^ in[46]); 
    assign layer_0[3677] = in[8]; 
    assign layer_0[3678] = ~(in[181] | in[164]); 
    assign layer_0[3679] = in[236] | in[158]; 
    assign layer_0[3680] = ~(in[22] | in[154]); 
    assign layer_0[3681] = in[248] | in[110]; 
    assign layer_0[3682] = in[43] ^ in[106]; 
    assign layer_0[3683] = ~in[126] | (in[126] & in[249]); 
    assign layer_0[3684] = in[124] ^ in[106]; 
    assign layer_0[3685] = ~(in[181] ^ in[199]); 
    assign layer_0[3686] = ~(in[133] ^ in[131]); 
    assign layer_0[3687] = in[78]; 
    assign layer_0[3688] = ~in[164] | (in[70] & in[164]); 
    assign layer_0[3689] = in[119] & in[246]; 
    assign layer_0[3690] = in[213]; 
    assign layer_0[3691] = ~(in[95] ^ in[153]); 
    assign layer_0[3692] = in[60] & ~in[136]; 
    assign layer_0[3693] = ~in[44] | (in[41] & in[44]); 
    assign layer_0[3694] = ~(in[197] & in[183]); 
    assign layer_0[3695] = ~(in[195] | in[187]); 
    assign layer_0[3696] = ~in[57]; 
    assign layer_0[3697] = ~(in[233] ^ in[202]); 
    assign layer_0[3698] = ~in[75] | (in[217] & in[75]); 
    assign layer_0[3699] = ~(in[187] ^ in[189]); 
    assign layer_0[3700] = in[5] ^ in[7]; 
    assign layer_0[3701] = ~in[47]; 
    assign layer_0[3702] = in[91] & ~in[27]; 
    assign layer_0[3703] = in[26] | in[9]; 
    assign layer_0[3704] = in[189] | in[89]; 
    assign layer_0[3705] = ~in[97] | (in[93] & in[97]); 
    assign layer_0[3706] = in[140] | in[184]; 
    assign layer_0[3707] = in[63] | in[10]; 
    assign layer_0[3708] = ~(in[139] ^ in[79]); 
    assign layer_0[3709] = ~(in[236] ^ in[212]); 
    assign layer_0[3710] = in[120]; 
    assign layer_0[3711] = ~in[132] | (in[82] & in[132]); 
    assign layer_0[3712] = ~(in[81] | in[103]); 
    assign layer_0[3713] = in[90] & ~in[233]; 
    assign layer_0[3714] = in[63] ^ in[28]; 
    assign layer_0[3715] = in[164] | in[135]; 
    assign layer_0[3716] = in[228] ^ in[79]; 
    assign layer_0[3717] = ~(in[241] ^ in[245]); 
    assign layer_0[3718] = ~(in[113] ^ in[110]); 
    assign layer_0[3719] = ~(in[82] ^ in[151]); 
    assign layer_0[3720] = ~(in[85] ^ in[7]); 
    assign layer_0[3721] = ~in[73] | (in[73] & in[135]); 
    assign layer_0[3722] = ~in[167] | (in[196] & in[167]); 
    assign layer_0[3723] = in[180] ^ in[245]; 
    assign layer_0[3724] = ~in[88] | (in[88] & in[136]); 
    assign layer_0[3725] = ~(in[196] | in[211]); 
    assign layer_0[3726] = in[131] | in[133]; 
    assign layer_0[3727] = ~in[104] | (in[67] & in[104]); 
    assign layer_0[3728] = in[88] ^ in[50]; 
    assign layer_0[3729] = ~in[221]; 
    assign layer_0[3730] = in[91] ^ in[89]; 
    assign layer_0[3731] = ~(in[107] ^ in[149]); 
    assign layer_0[3732] = in[57] & ~in[157]; 
    assign layer_0[3733] = ~(in[140] & in[147]); 
    assign layer_0[3734] = in[125] ^ in[123]; 
    assign layer_0[3735] = ~(in[76] & in[109]); 
    assign layer_0[3736] = in[133] ^ in[163]; 
    assign layer_0[3737] = ~(in[74] | in[252]); 
    assign layer_0[3738] = in[103]; 
    assign layer_0[3739] = ~(in[178] | in[235]); 
    assign layer_0[3740] = in[120] ^ in[166]; 
    assign layer_0[3741] = in[103] & ~in[84]; 
    assign layer_0[3742] = in[58] | in[88]; 
    assign layer_0[3743] = ~(in[230] | in[199]); 
    assign layer_0[3744] = ~(in[248] | in[202]); 
    assign layer_0[3745] = in[233] ^ in[242]; 
    assign layer_0[3746] = in[69] & ~in[117]; 
    assign layer_0[3747] = ~(in[52] | in[24]); 
    assign layer_0[3748] = ~in[220]; 
    assign layer_0[3749] = ~(in[245] ^ in[214]); 
    assign layer_0[3750] = ~(in[76] ^ in[107]); 
    assign layer_0[3751] = ~(in[226] ^ in[181]); 
    assign layer_0[3752] = ~(in[10] | in[71]); 
    assign layer_0[3753] = in[80] ^ in[242]; 
    assign layer_0[3754] = in[152] | in[212]; 
    assign layer_0[3755] = in[22] ^ in[56]; 
    assign layer_0[3756] = ~in[157]; 
    assign layer_0[3757] = in[92] ^ in[51]; 
    assign layer_0[3758] = ~in[184] | (in[184] & in[126]); 
    assign layer_0[3759] = in[115] ^ in[101]; 
    assign layer_0[3760] = in[169] & in[78]; 
    assign layer_0[3761] = ~in[249]; 
    assign layer_0[3762] = in[180] ^ in[178]; 
    assign layer_0[3763] = in[168] | in[107]; 
    assign layer_0[3764] = ~(in[39] | in[213]); 
    assign layer_0[3765] = ~(in[198] | in[206]); 
    assign layer_0[3766] = ~(in[81] | in[73]); 
    assign layer_0[3767] = ~in[246] | (in[246] & in[25]); 
    assign layer_0[3768] = ~(in[108] ^ in[139]); 
    assign layer_0[3769] = ~in[184] | (in[40] & in[184]); 
    assign layer_0[3770] = in[199] ^ in[92]; 
    assign layer_0[3771] = in[29] ^ in[62]; 
    assign layer_0[3772] = ~(in[247] ^ in[241]); 
    assign layer_0[3773] = in[200] ^ in[167]; 
    assign layer_0[3774] = ~(in[220] ^ in[111]); 
    assign layer_0[3775] = in[166] ^ in[121]; 
    assign layer_0[3776] = ~(in[77] | in[214]); 
    assign layer_0[3777] = ~(in[251] ^ in[219]); 
    assign layer_0[3778] = ~in[131] | (in[131] & in[219]); 
    assign layer_0[3779] = in[74] ^ in[119]; 
    assign layer_0[3780] = ~(in[245] ^ in[212]); 
    assign layer_0[3781] = in[235] ^ in[218]; 
    assign layer_0[3782] = ~(in[41] | in[44]); 
    assign layer_0[3783] = ~(in[166] ^ in[164]); 
    assign layer_0[3784] = in[53] ^ in[21]; 
    assign layer_0[3785] = in[140] ^ in[171]; 
    assign layer_0[3786] = ~(in[142] | in[250]); 
    assign layer_0[3787] = in[164] | in[125]; 
    assign layer_0[3788] = in[51] | in[149]; 
    assign layer_0[3789] = in[102] ^ in[23]; 
    assign layer_0[3790] = ~(in[184] & in[51]); 
    assign layer_0[3791] = ~in[66]; 
    assign layer_0[3792] = in[74] | in[72]; 
    assign layer_0[3793] = in[125] | in[122]; 
    assign layer_0[3794] = in[43] | in[180]; 
    assign layer_0[3795] = in[51] ^ in[155]; 
    assign layer_0[3796] = in[90] | in[78]; 
    assign layer_0[3797] = ~(in[234] ^ in[216]); 
    assign layer_0[3798] = ~(in[203] ^ in[38]); 
    assign layer_0[3799] = in[41] & ~in[39]; 
    assign layer_0[3800] = in[56] & ~in[210]; 
    assign layer_0[3801] = in[104] & ~in[133]; 
    assign layer_0[3802] = ~(in[72] | in[93]); 
    assign layer_0[3803] = ~(in[78] | in[51]); 
    assign layer_0[3804] = ~(in[27] | in[150]); 
    assign layer_0[3805] = in[91]; 
    assign layer_0[3806] = in[168] & ~in[163]; 
    assign layer_0[3807] = ~(in[125] | in[170]); 
    assign layer_0[3808] = in[135] | in[228]; 
    assign layer_0[3809] = in[53] ^ in[99]; 
    assign layer_0[3810] = ~in[165]; 
    assign layer_0[3811] = ~(in[108] ^ in[110]); 
    assign layer_0[3812] = in[41] ^ in[29]; 
    assign layer_0[3813] = in[205] | in[25]; 
    assign layer_0[3814] = in[72] & ~in[108]; 
    assign layer_0[3815] = ~(in[95] | in[161]); 
    assign layer_0[3816] = ~(in[22] | in[156]); 
    assign layer_0[3817] = ~(in[146] | in[166]); 
    assign layer_0[3818] = ~(in[27] | in[213]); 
    assign layer_0[3819] = ~(in[149] | in[95]); 
    assign layer_0[3820] = ~(in[73] | in[77]); 
    assign layer_0[3821] = ~(in[124] | in[90]); 
    assign layer_0[3822] = in[23] ^ in[186]; 
    assign layer_0[3823] = in[102] ^ in[170]; 
    assign layer_0[3824] = ~in[105] | (in[139] & in[105]); 
    assign layer_0[3825] = ~(in[134] | in[193]); 
    assign layer_0[3826] = ~in[142] | (in[229] & in[142]); 
    assign layer_0[3827] = in[119] ^ in[150]; 
    assign layer_0[3828] = ~(in[50] ^ in[210]); 
    assign layer_0[3829] = in[120] & ~in[107]; 
    assign layer_0[3830] = in[100] | in[149]; 
    assign layer_0[3831] = in[181] ^ in[179]; 
    assign layer_0[3832] = ~in[35]; 
    assign layer_0[3833] = in[233] ^ in[188]; 
    assign layer_0[3834] = in[36] | in[107]; 
    assign layer_0[3835] = in[74] & in[42]; 
    assign layer_0[3836] = ~(in[59] | in[56]); 
    assign layer_0[3837] = in[105] ^ in[125]; 
    assign layer_0[3838] = ~(in[248] | in[106]); 
    assign layer_0[3839] = in[136] | in[6]; 
    assign layer_0[3840] = in[137]; 
    assign layer_0[3841] = ~in[167] | (in[110] & in[167]); 
    assign layer_0[3842] = in[164] | in[168]; 
    assign layer_0[3843] = ~(in[180] | in[162]); 
    assign layer_0[3844] = in[132] ^ in[146]; 
    assign layer_0[3845] = ~(in[227] ^ in[72]); 
    assign layer_0[3846] = ~(in[93] | in[80]); 
    assign layer_0[3847] = ~(in[143] | in[35]); 
    assign layer_0[3848] = ~(in[126] | in[196]); 
    assign layer_0[3849] = ~(in[155] | in[155]); 
    assign layer_0[3850] = ~in[202] | (in[202] & in[131]); 
    assign layer_0[3851] = ~in[170]; 
    assign layer_0[3852] = ~(in[181] ^ in[229]); 
    assign layer_0[3853] = in[213]; 
    assign layer_0[3854] = ~(in[58] ^ in[89]); 
    assign layer_0[3855] = ~(in[241] | in[173]); 
    assign layer_0[3856] = in[156] | in[199]; 
    assign layer_0[3857] = ~(in[119] ^ in[149]); 
    assign layer_0[3858] = in[58] ^ in[90]; 
    assign layer_0[3859] = in[157] | in[243]; 
    assign layer_0[3860] = in[182] & ~in[236]; 
    assign layer_0[3861] = ~(in[199] ^ in[136]); 
    assign layer_0[3862] = in[79] | in[235]; 
    assign layer_0[3863] = in[214] & ~in[89]; 
    assign layer_0[3864] = ~(in[149] | in[124]); 
    assign layer_0[3865] = in[104] & ~in[92]; 
    assign layer_0[3866] = in[152] & ~in[10]; 
    assign layer_0[3867] = in[123]; 
    assign layer_0[3868] = in[170] & ~in[104]; 
    assign layer_0[3869] = ~(in[104] | in[231]); 
    assign layer_0[3870] = in[229] | in[231]; 
    assign layer_0[3871] = ~in[155] | (in[221] & in[155]); 
    assign layer_0[3872] = in[189] | in[219]; 
    assign layer_0[3873] = ~(in[202] | in[233]); 
    assign layer_0[3874] = ~in[215]; 
    assign layer_0[3875] = ~(in[83] | in[178]); 
    assign layer_0[3876] = ~(in[44] ^ in[186]); 
    assign layer_0[3877] = ~(in[10] ^ in[59]); 
    assign layer_0[3878] = ~(in[22] ^ in[162]); 
    assign layer_0[3879] = in[185] ^ in[103]; 
    assign layer_0[3880] = ~(in[206] | in[120]); 
    assign layer_0[3881] = in[227]; 
    assign layer_0[3882] = ~in[86]; 
    assign layer_0[3883] = ~(in[243] ^ in[155]); 
    assign layer_0[3884] = in[36] | in[25]; 
    assign layer_0[3885] = in[41] & ~in[109]; 
    assign layer_0[3886] = ~(in[11] | in[28]); 
    assign layer_0[3887] = in[170] ^ in[59]; 
    assign layer_0[3888] = in[152] ^ in[177]; 
    assign layer_0[3889] = in[181] & ~in[6]; 
    assign layer_0[3890] = ~in[153] | (in[153] & in[164]); 
    assign layer_0[3891] = ~(in[237] | in[191]); 
    assign layer_0[3892] = ~(in[132] ^ in[196]); 
    assign layer_0[3893] = ~(in[232] ^ in[185]); 
    assign layer_0[3894] = in[116] ^ in[102]; 
    assign layer_0[3895] = in[163] | in[131]; 
    assign layer_0[3896] = in[233] | in[180]; 
    assign layer_0[3897] = ~in[234] | (in[234] & in[121]); 
    assign layer_0[3898] = in[104] | in[25]; 
    assign layer_0[3899] = ~(in[163] | in[130]); 
    assign layer_0[3900] = ~(in[193] | in[179]); 
    assign layer_0[3901] = in[46]; 
    assign layer_0[3902] = in[102] ^ in[243]; 
    assign layer_0[3903] = ~(in[199] ^ in[44]); 
    assign layer_0[3904] = in[86] ^ in[67]; 
    assign layer_0[3905] = ~in[221]; 
    assign layer_0[3906] = ~in[70] | (in[70] & in[83]); 
    assign layer_0[3907] = ~in[53]; 
    assign layer_0[3908] = ~in[87] | (in[251] & in[87]); 
    assign layer_0[3909] = ~(in[133] ^ in[75]); 
    assign layer_0[3910] = in[86] & ~in[135]; 
    assign layer_0[3911] = ~(in[248] ^ in[185]); 
    assign layer_0[3912] = in[229] & ~in[219]; 
    assign layer_0[3913] = ~in[126] | (in[126] & in[135]); 
    assign layer_0[3914] = ~(in[131] | in[227]); 
    assign layer_0[3915] = ~(in[118] | in[148]); 
    assign layer_0[3916] = ~(in[110] ^ in[108]); 
    assign layer_0[3917] = ~(in[115] ^ in[117]); 
    assign layer_0[3918] = in[68]; 
    assign layer_0[3919] = in[182]; 
    assign layer_0[3920] = in[104] & ~in[107]; 
    assign layer_0[3921] = in[195] ^ in[143]; 
    assign layer_0[3922] = ~in[103] | (in[103] & in[69]); 
    assign layer_0[3923] = ~in[154] | (in[141] & in[154]); 
    assign layer_0[3924] = in[72] & in[58]; 
    assign layer_0[3925] = in[35] | in[176]; 
    assign layer_0[3926] = in[19]; 
    assign layer_0[3927] = in[180] ^ in[105]; 
    assign layer_0[3928] = in[39] ^ in[8]; 
    assign layer_0[3929] = ~(in[52] ^ in[82]); 
    assign layer_0[3930] = in[130] ^ in[39]; 
    assign layer_0[3931] = in[217] & ~in[83]; 
    assign layer_0[3932] = ~(in[132] | in[130]); 
    assign layer_0[3933] = in[69] ^ in[23]; 
    assign layer_0[3934] = in[76]; 
    assign layer_0[3935] = ~(in[89] | in[123]); 
    assign layer_0[3936] = in[72] ^ in[195]; 
    assign layer_0[3937] = ~in[215] | (in[215] & in[229]); 
    assign layer_0[3938] = in[248] | in[118]; 
    assign layer_0[3939] = ~(in[89] ^ in[104]); 
    assign layer_0[3940] = in[226] | in[209]; 
    assign layer_0[3941] = ~in[130]; 
    assign layer_0[3942] = in[103]; 
    assign layer_0[3943] = in[102]; 
    assign layer_0[3944] = ~in[85] | (in[85] & in[148]); 
    assign layer_0[3945] = ~(in[114] ^ in[101]); 
    assign layer_0[3946] = in[150] | in[82]; 
    assign layer_0[3947] = ~(in[76] | in[215]); 
    assign layer_0[3948] = in[73] | in[41]; 
    assign layer_0[3949] = ~in[217] | (in[217] & in[171]); 
    assign layer_0[3950] = ~in[85]; 
    assign layer_0[3951] = ~in[10] | (in[10] & in[228]); 
    assign layer_0[3952] = ~(in[69] ^ in[102]); 
    assign layer_0[3953] = ~(in[74] & in[69]); 
    assign layer_0[3954] = in[250] | in[108]; 
    assign layer_0[3955] = ~(in[204] ^ in[201]); 
    assign layer_0[3956] = in[230] ^ in[183]; 
    assign layer_0[3957] = in[101] & ~in[214]; 
    assign layer_0[3958] = ~(in[124] ^ in[166]); 
    assign layer_0[3959] = ~in[170] | (in[170] & in[204]); 
    assign layer_0[3960] = in[163]; 
    assign layer_0[3961] = in[115] ^ in[117]; 
    assign layer_0[3962] = ~in[218] | (in[218] & in[125]); 
    assign layer_0[3963] = ~(in[156] ^ in[137]); 
    assign layer_0[3964] = in[87] ^ in[116]; 
    assign layer_0[3965] = ~(in[71] ^ in[38]); 
    assign layer_0[3966] = ~(in[126] | in[214]); 
    assign layer_0[3967] = ~in[71] | (in[71] & in[52]); 
    assign layer_0[3968] = ~in[116] | (in[116] & in[9]); 
    assign layer_0[3969] = ~in[67]; 
    assign layer_0[3970] = in[151] ^ in[104]; 
    assign layer_0[3971] = in[212] ^ in[94]; 
    assign layer_0[3972] = ~(in[76] | in[107]); 
    assign layer_0[3973] = ~in[136] | (in[76] & in[136]); 
    assign layer_0[3974] = ~(in[55] & in[70]); 
    assign layer_0[3975] = ~(in[199] ^ in[246]); 
    assign layer_0[3976] = ~(in[183] ^ in[122]); 
    assign layer_0[3977] = ~(in[185] ^ in[242]); 
    assign layer_0[3978] = ~in[182] | (in[182] & in[78]); 
    assign layer_0[3979] = ~(in[36] | in[21]); 
    assign layer_0[3980] = in[93] | in[228]; 
    assign layer_0[3981] = in[167] & ~in[20]; 
    assign layer_0[3982] = in[63] | in[139]; 
    assign layer_0[3983] = ~(in[83] ^ in[69]); 
    assign layer_0[3984] = ~in[178] | (in[178] & in[232]); 
    assign layer_0[3985] = in[37] | in[171]; 
    assign layer_0[3986] = in[121] ^ in[131]; 
    assign layer_0[3987] = in[218] ^ in[81]; 
    assign layer_0[3988] = ~(in[158] | in[62]); 
    assign layer_0[3989] = in[82] | in[40]; 
    assign layer_0[3990] = in[21] ^ in[143]; 
    assign layer_0[3991] = in[52] ^ in[81]; 
    assign layer_0[3992] = ~in[138] | (in[41] & in[138]); 
    assign layer_0[3993] = ~(in[102] ^ in[70]); 
    assign layer_0[3994] = ~(in[183] ^ in[181]); 
    assign layer_0[3995] = ~(in[60] ^ in[91]); 
    assign layer_0[3996] = in[218] ^ in[183]; 
    assign layer_0[3997] = ~(in[107] ^ in[125]); 
    assign layer_0[3998] = in[121] ^ in[140]; 
    assign layer_0[3999] = in[91] ^ in[93]; 
    // Layer 1 ============================================================
    assign out[0] = layer_0[1562] & layer_0[2267]; 
    assign out[1] = layer_0[3041] ^ layer_0[2261]; 
    assign out[2] = layer_0[3485] & layer_0[1315]; 
    assign out[3] = layer_0[2208] ^ layer_0[1920]; 
    assign out[4] = ~layer_0[372]; 
    assign out[5] = ~layer_0[3332] | (layer_0[2259] & layer_0[3332]); 
    assign out[6] = layer_0[3377] & ~layer_0[349]; 
    assign out[7] = ~(layer_0[3946] | layer_0[358]); 
    assign out[8] = layer_0[3973] & ~layer_0[3263]; 
    assign out[9] = layer_0[2007] & layer_0[3393]; 
    assign out[10] = ~layer_0[1561] | (layer_0[1561] & layer_0[1419]); 
    assign out[11] = ~layer_0[2858]; 
    assign out[12] = ~layer_0[1166]; 
    assign out[13] = layer_0[1488] ^ layer_0[2803]; 
    assign out[14] = ~(layer_0[3528] & layer_0[2541]); 
    assign out[15] = ~layer_0[1105]; 
    assign out[16] = ~layer_0[3033]; 
    assign out[17] = ~layer_0[3193]; 
    assign out[18] = layer_0[2774] & ~layer_0[2228]; 
    assign out[19] = ~layer_0[2453]; 
    assign out[20] = layer_0[2079] & ~layer_0[386]; 
    assign out[21] = layer_0[1740] ^ layer_0[1670]; 
    assign out[22] = layer_0[2515] & ~layer_0[3598]; 
    assign out[23] = ~(layer_0[2178] ^ layer_0[2894]); 
    assign out[24] = layer_0[3272] & ~layer_0[2764]; 
    assign out[25] = layer_0[1191] & ~layer_0[1758]; 
    assign out[26] = ~layer_0[2205]; 
    assign out[27] = layer_0[3622] & ~layer_0[1926]; 
    assign out[28] = ~layer_0[2390]; 
    assign out[29] = layer_0[196] & ~layer_0[534]; 
    assign out[30] = layer_0[262] ^ layer_0[1149]; 
    assign out[31] = layer_0[548] ^ layer_0[3966]; 
    assign out[32] = layer_0[1007] ^ layer_0[2899]; 
    assign out[33] = layer_0[1053] & ~layer_0[521]; 
    assign out[34] = layer_0[868] & ~layer_0[1737]; 
    assign out[35] = ~(layer_0[3688] & layer_0[1333]); 
    assign out[36] = ~layer_0[3823]; 
    assign out[37] = layer_0[2901]; 
    assign out[38] = ~layer_0[3652] | (layer_0[3652] & layer_0[2040]); 
    assign out[39] = ~(layer_0[134] ^ layer_0[304]); 
    assign out[40] = layer_0[3731]; 
    assign out[41] = layer_0[3209] ^ layer_0[3034]; 
    assign out[42] = ~layer_0[1129]; 
    assign out[43] = layer_0[2006] & ~layer_0[2189]; 
    assign out[44] = ~layer_0[1087]; 
    assign out[45] = layer_0[776] ^ layer_0[3783]; 
    assign out[46] = layer_0[1701] | layer_0[952]; 
    assign out[47] = layer_0[708] ^ layer_0[1411]; 
    assign out[48] = layer_0[3399] ^ layer_0[3241]; 
    assign out[49] = ~layer_0[405] | (layer_0[405] & layer_0[2986]); 
    assign out[50] = layer_0[1568] & layer_0[2989]; 
    assign out[51] = layer_0[3146]; 
    assign out[52] = layer_0[3196] & ~layer_0[330]; 
    assign out[53] = layer_0[263] & ~layer_0[1377]; 
    assign out[54] = layer_0[435] & layer_0[3890]; 
    assign out[55] = layer_0[391] ^ layer_0[2913]; 
    assign out[56] = ~(layer_0[3242] ^ layer_0[324]); 
    assign out[57] = ~(layer_0[549] & layer_0[3671]); 
    assign out[58] = ~(layer_0[371] ^ layer_0[362]); 
    assign out[59] = layer_0[2524] & ~layer_0[1407]; 
    assign out[60] = layer_0[2791]; 
    assign out[61] = layer_0[1291]; 
    assign out[62] = ~layer_0[2244]; 
    assign out[63] = layer_0[1026] & ~layer_0[2043]; 
    assign out[64] = ~layer_0[1300]; 
    assign out[65] = layer_0[75] ^ layer_0[3602]; 
    assign out[66] = layer_0[566] ^ layer_0[1691]; 
    assign out[67] = ~(layer_0[51] | layer_0[89]); 
    assign out[68] = layer_0[1653] ^ layer_0[2998]; 
    assign out[69] = layer_0[1543] ^ layer_0[676]; 
    assign out[70] = layer_0[1201] ^ layer_0[1906]; 
    assign out[71] = layer_0[1243]; 
    assign out[72] = layer_0[3268] ^ layer_0[1841]; 
    assign out[73] = layer_0[2261] & layer_0[3976]; 
    assign out[74] = layer_0[1433]; 
    assign out[75] = ~(layer_0[2437] & layer_0[2406]); 
    assign out[76] = layer_0[2549] & layer_0[2315]; 
    assign out[77] = layer_0[1019] & ~layer_0[3035]; 
    assign out[78] = ~(layer_0[1151] | layer_0[3351]); 
    assign out[79] = layer_0[1615] & ~layer_0[490]; 
    assign out[80] = layer_0[562]; 
    assign out[81] = ~layer_0[1414]; 
    assign out[82] = ~(layer_0[3415] ^ layer_0[2949]); 
    assign out[83] = ~layer_0[588]; 
    assign out[84] = layer_0[1911] & layer_0[3140]; 
    assign out[85] = ~(layer_0[280] | layer_0[7]); 
    assign out[86] = layer_0[518]; 
    assign out[87] = layer_0[3973]; 
    assign out[88] = ~(layer_0[211] | layer_0[1452]); 
    assign out[89] = layer_0[3591]; 
    assign out[90] = ~(layer_0[224] ^ layer_0[846]); 
    assign out[91] = layer_0[1191]; 
    assign out[92] = layer_0[3435]; 
    assign out[93] = layer_0[3371] & ~layer_0[2465]; 
    assign out[94] = layer_0[1728]; 
    assign out[95] = ~layer_0[462]; 
    assign out[96] = layer_0[306] ^ layer_0[1721]; 
    assign out[97] = ~(layer_0[2983] | layer_0[2992]); 
    assign out[98] = ~layer_0[311] | (layer_0[311] & layer_0[3880]); 
    assign out[99] = ~(layer_0[1798] ^ layer_0[903]); 
    assign out[100] = ~(layer_0[1865] ^ layer_0[3758]); 
    assign out[101] = layer_0[2061]; 
    assign out[102] = ~(layer_0[1233] ^ layer_0[325]); 
    assign out[103] = layer_0[990] & ~layer_0[3551]; 
    assign out[104] = layer_0[1231]; 
    assign out[105] = ~(layer_0[102] ^ layer_0[3995]); 
    assign out[106] = ~(layer_0[1024] | layer_0[431]); 
    assign out[107] = ~layer_0[1833]; 
    assign out[108] = layer_0[3087]; 
    assign out[109] = ~layer_0[3389] | (layer_0[3389] & layer_0[608]); 
    assign out[110] = layer_0[1775] ^ layer_0[1978]; 
    assign out[111] = ~(layer_0[3683] ^ layer_0[1666]); 
    assign out[112] = layer_0[2696] & layer_0[1795]; 
    assign out[113] = layer_0[3516] & layer_0[1842]; 
    assign out[114] = ~layer_0[2129]; 
    assign out[115] = layer_0[1979]; 
    assign out[116] = layer_0[2381] & ~layer_0[722]; 
    assign out[117] = layer_0[1732] & ~layer_0[922]; 
    assign out[118] = ~(layer_0[249] ^ layer_0[1155]); 
    assign out[119] = layer_0[1573]; 
    assign out[120] = ~(layer_0[1809] | layer_0[112]); 
    assign out[121] = ~(layer_0[1254] ^ layer_0[3761]); 
    assign out[122] = ~layer_0[2594] | (layer_0[2105] & layer_0[2594]); 
    assign out[123] = ~layer_0[3143]; 
    assign out[124] = layer_0[799] & ~layer_0[1379]; 
    assign out[125] = layer_0[3333] ^ layer_0[2746]; 
    assign out[126] = ~layer_0[1874] | (layer_0[3434] & layer_0[1874]); 
    assign out[127] = layer_0[2590] & layer_0[3368]; 
    assign out[128] = ~(layer_0[2574] | layer_0[1418]); 
    assign out[129] = ~layer_0[3749]; 
    assign out[130] = layer_0[1702]; 
    assign out[131] = layer_0[1476]; 
    assign out[132] = layer_0[796] ^ layer_0[1423]; 
    assign out[133] = ~(layer_0[610] | layer_0[1202]); 
    assign out[134] = layer_0[2026] ^ layer_0[3092]; 
    assign out[135] = ~layer_0[2383] | (layer_0[2383] & layer_0[1729]); 
    assign out[136] = layer_0[1870]; 
    assign out[137] = layer_0[623] & layer_0[3309]; 
    assign out[138] = ~layer_0[172] | (layer_0[2278] & layer_0[172]); 
    assign out[139] = layer_0[1011] ^ layer_0[1413]; 
    assign out[140] = ~(layer_0[1247] & layer_0[2617]); 
    assign out[141] = layer_0[2966]; 
    assign out[142] = layer_0[3038] & ~layer_0[1827]; 
    assign out[143] = ~(layer_0[707] ^ layer_0[1477]); 
    assign out[144] = layer_0[2374] & layer_0[3961]; 
    assign out[145] = ~(layer_0[165] | layer_0[2919]); 
    assign out[146] = ~(layer_0[1783] ^ layer_0[2168]); 
    assign out[147] = ~layer_0[1539] | (layer_0[1539] & layer_0[3259]); 
    assign out[148] = ~layer_0[2857]; 
    assign out[149] = ~layer_0[2454] | (layer_0[2454] & layer_0[904]); 
    assign out[150] = layer_0[1344] ^ layer_0[316]; 
    assign out[151] = layer_0[3634] ^ layer_0[84]; 
    assign out[152] = ~(layer_0[965] ^ layer_0[2368]); 
    assign out[153] = layer_0[1292] & ~layer_0[2246]; 
    assign out[154] = ~layer_0[1977]; 
    assign out[155] = layer_0[2128] & ~layer_0[2133]; 
    assign out[156] = layer_0[1471]; 
    assign out[157] = ~(layer_0[82] ^ layer_0[879]); 
    assign out[158] = layer_0[2230] & layer_0[3414]; 
    assign out[159] = ~(layer_0[620] & layer_0[2634]); 
    assign out[160] = layer_0[116] ^ layer_0[877]; 
    assign out[161] = ~layer_0[1710]; 
    assign out[162] = layer_0[1952] ^ layer_0[969]; 
    assign out[163] = layer_0[1355] ^ layer_0[3943]; 
    assign out[164] = ~layer_0[3743]; 
    assign out[165] = layer_0[1844]; 
    assign out[166] = layer_0[3379] & ~layer_0[446]; 
    assign out[167] = ~layer_0[1058] | (layer_0[2103] & layer_0[1058]); 
    assign out[168] = layer_0[2732]; 
    assign out[169] = ~(layer_0[250] | layer_0[443]); 
    assign out[170] = layer_0[2293] & ~layer_0[921]; 
    assign out[171] = layer_0[393]; 
    assign out[172] = ~layer_0[3879]; 
    assign out[173] = ~(layer_0[717] ^ layer_0[2315]); 
    assign out[174] = ~layer_0[3827]; 
    assign out[175] = ~(layer_0[3219] ^ layer_0[3597]); 
    assign out[176] = layer_0[3545] & layer_0[2323]; 
    assign out[177] = ~layer_0[179]; 
    assign out[178] = ~layer_0[537]; 
    assign out[179] = ~layer_0[1741]; 
    assign out[180] = ~layer_0[2225] | (layer_0[2225] & layer_0[1724]); 
    assign out[181] = ~(layer_0[2948] | layer_0[750]); 
    assign out[182] = ~layer_0[636]; 
    assign out[183] = ~(layer_0[1121] ^ layer_0[175]); 
    assign out[184] = layer_0[1122] | layer_0[1965]; 
    assign out[185] = layer_0[2572] ^ layer_0[1776]; 
    assign out[186] = ~(layer_0[3017] | layer_0[3913]); 
    assign out[187] = ~(layer_0[1891] | layer_0[2455]); 
    assign out[188] = layer_0[1779] ^ layer_0[1088]; 
    assign out[189] = ~(layer_0[349] | layer_0[2467]); 
    assign out[190] = layer_0[1972] ^ layer_0[2741]; 
    assign out[191] = layer_0[417] ^ layer_0[3510]; 
    assign out[192] = ~(layer_0[1968] | layer_0[351]); 
    assign out[193] = ~(layer_0[931] | layer_0[2759]); 
    assign out[194] = layer_0[2143] & layer_0[536]; 
    assign out[195] = ~layer_0[571] | (layer_0[632] & layer_0[571]); 
    assign out[196] = layer_0[1910]; 
    assign out[197] = layer_0[221] ^ layer_0[3232]; 
    assign out[198] = ~(layer_0[38] ^ layer_0[245]); 
    assign out[199] = layer_0[1204] ^ layer_0[270]; 
    assign out[200] = layer_0[3637] & ~layer_0[3360]; 
    assign out[201] = layer_0[1187]; 
    assign out[202] = layer_0[3243] & ~layer_0[2314]; 
    assign out[203] = ~layer_0[1706]; 
    assign out[204] = layer_0[268]; 
    assign out[205] = ~layer_0[3413]; 
    assign out[206] = layer_0[2659] & layer_0[1842]; 
    assign out[207] = ~(layer_0[2411] | layer_0[768]); 
    assign out[208] = ~layer_0[386]; 
    assign out[209] = ~layer_0[2763]; 
    assign out[210] = layer_0[2704]; 
    assign out[211] = ~(layer_0[1039] ^ layer_0[401]); 
    assign out[212] = ~(layer_0[3482] | layer_0[2762]); 
    assign out[213] = layer_0[2443]; 
    assign out[214] = ~(layer_0[2961] ^ layer_0[482]); 
    assign out[215] = layer_0[1329]; 
    assign out[216] = ~(layer_0[2197] ^ layer_0[1252]); 
    assign out[217] = ~layer_0[458] | (layer_0[458] & layer_0[3546]); 
    assign out[218] = layer_0[2365] ^ layer_0[3354]; 
    assign out[219] = layer_0[3010] & ~layer_0[3848]; 
    assign out[220] = ~(layer_0[1580] | layer_0[1836]); 
    assign out[221] = ~layer_0[3666]; 
    assign out[222] = ~(layer_0[3203] ^ layer_0[1950]); 
    assign out[223] = layer_0[3556] | layer_0[3661]; 
    assign out[224] = layer_0[1575] & ~layer_0[3202]; 
    assign out[225] = ~(layer_0[26] ^ layer_0[3088]); 
    assign out[226] = ~(layer_0[2866] | layer_0[2573]); 
    assign out[227] = layer_0[427]; 
    assign out[228] = ~(layer_0[438] ^ layer_0[2197]); 
    assign out[229] = layer_0[781]; 
    assign out[230] = layer_0[2094] & ~layer_0[1072]; 
    assign out[231] = layer_0[3656] ^ layer_0[1838]; 
    assign out[232] = ~layer_0[1441]; 
    assign out[233] = layer_0[791] & layer_0[1411]; 
    assign out[234] = layer_0[583]; 
    assign out[235] = ~layer_0[2456] | (layer_0[2456] & layer_0[303]); 
    assign out[236] = ~(layer_0[1985] ^ layer_0[3457]); 
    assign out[237] = ~layer_0[383]; 
    assign out[238] = layer_0[484] ^ layer_0[2090]; 
    assign out[239] = layer_0[1757] ^ layer_0[3769]; 
    assign out[240] = layer_0[1219] ^ layer_0[2212]; 
    assign out[241] = layer_0[399] & ~layer_0[2313]; 
    assign out[242] = ~(layer_0[1893] ^ layer_0[1595]); 
    assign out[243] = ~layer_0[3623]; 
    assign out[244] = ~(layer_0[3021] ^ layer_0[1168]); 
    assign out[245] = ~(layer_0[811] ^ layer_0[3912]); 
    assign out[246] = ~(layer_0[2931] ^ layer_0[2220]); 
    assign out[247] = ~(layer_0[3900] ^ layer_0[2814]); 
    assign out[248] = layer_0[2625]; 
    assign out[249] = layer_0[847] ^ layer_0[3240]; 
    assign out[250] = ~layer_0[2693] | (layer_0[2693] & layer_0[2533]); 
    assign out[251] = ~(layer_0[340] ^ layer_0[1159]); 
    assign out[252] = ~(layer_0[2753] | layer_0[1672]); 
    assign out[253] = ~layer_0[871] | (layer_0[871] & layer_0[1564]); 
    assign out[254] = ~(layer_0[2882] & layer_0[269]); 
    assign out[255] = ~layer_0[1638] | (layer_0[1638] & layer_0[93]); 
    assign out[256] = layer_0[2957]; 
    assign out[257] = ~(layer_0[3875] ^ layer_0[227]); 
    assign out[258] = layer_0[979] | layer_0[3354]; 
    assign out[259] = ~layer_0[1604]; 
    assign out[260] = layer_0[508] ^ layer_0[138]; 
    assign out[261] = layer_0[1681] & layer_0[1709]; 
    assign out[262] = ~(layer_0[2745] ^ layer_0[1959]); 
    assign out[263] = ~layer_0[3032]; 
    assign out[264] = layer_0[17] ^ layer_0[1496]; 
    assign out[265] = ~(layer_0[756] ^ layer_0[1602]); 
    assign out[266] = ~layer_0[2060] | (layer_0[2060] & layer_0[96]); 
    assign out[267] = layer_0[3474]; 
    assign out[268] = ~(layer_0[3822] | layer_0[1363]); 
    assign out[269] = layer_0[3770]; 
    assign out[270] = layer_0[180] ^ layer_0[3788]; 
    assign out[271] = layer_0[390] & layer_0[1565]; 
    assign out[272] = layer_0[2518]; 
    assign out[273] = ~(layer_0[593] ^ layer_0[945]); 
    assign out[274] = layer_0[181] & ~layer_0[1280]; 
    assign out[275] = ~layer_0[523]; 
    assign out[276] = ~layer_0[40] | (layer_0[40] & layer_0[430]); 
    assign out[277] = ~(layer_0[2579] | layer_0[2210]); 
    assign out[278] = ~(layer_0[717] ^ layer_0[907]); 
    assign out[279] = layer_0[2413] & ~layer_0[1661]; 
    assign out[280] = layer_0[2641] ^ layer_0[2845]; 
    assign out[281] = ~(layer_0[2235] ^ layer_0[1499]); 
    assign out[282] = layer_0[3080] ^ layer_0[3554]; 
    assign out[283] = layer_0[1850]; 
    assign out[284] = ~layer_0[3392]; 
    assign out[285] = ~(layer_0[3011] ^ layer_0[2127]); 
    assign out[286] = ~(layer_0[1065] ^ layer_0[2175]); 
    assign out[287] = ~(layer_0[2812] & layer_0[3533]); 
    assign out[288] = layer_0[1364] & layer_0[3640]; 
    assign out[289] = layer_0[1351] & layer_0[2198]; 
    assign out[290] = ~(layer_0[3269] | layer_0[2761]); 
    assign out[291] = ~(layer_0[431] ^ layer_0[1115]); 
    assign out[292] = ~(layer_0[2274] | layer_0[4]); 
    assign out[293] = ~layer_0[3493]; 
    assign out[294] = layer_0[3119] & ~layer_0[3588]; 
    assign out[295] = ~(layer_0[1212] ^ layer_0[1894]); 
    assign out[296] = ~(layer_0[3462] ^ layer_0[3982]); 
    assign out[297] = layer_0[3768] | layer_0[544]; 
    assign out[298] = layer_0[865] & ~layer_0[317]; 
    assign out[299] = ~(layer_0[3483] | layer_0[951]); 
    assign out[300] = layer_0[2053] & ~layer_0[3004]; 
    assign out[301] = layer_0[2897] ^ layer_0[3834]; 
    assign out[302] = layer_0[744] & ~layer_0[3638]; 
    assign out[303] = layer_0[186] & layer_0[1617]; 
    assign out[304] = ~layer_0[625]; 
    assign out[305] = layer_0[1059] ^ layer_0[2355]; 
    assign out[306] = ~layer_0[3058]; 
    assign out[307] = layer_0[2216] & ~layer_0[1804]; 
    assign out[308] = layer_0[1745]; 
    assign out[309] = layer_0[3353]; 
    assign out[310] = layer_0[542] ^ layer_0[1685]; 
    assign out[311] = ~(layer_0[2548] | layer_0[964]); 
    assign out[312] = layer_0[3695] & ~layer_0[1584]; 
    assign out[313] = ~(layer_0[1782] ^ layer_0[278]); 
    assign out[314] = layer_0[1578] ^ layer_0[2029]; 
    assign out[315] = layer_0[3909]; 
    assign out[316] = ~(layer_0[2793] ^ layer_0[2142]); 
    assign out[317] = ~(layer_0[2880] ^ layer_0[3952]); 
    assign out[318] = layer_0[2349] & ~layer_0[1620]; 
    assign out[319] = ~(layer_0[580] ^ layer_0[1678]); 
    assign out[320] = ~layer_0[241]; 
    assign out[321] = ~(layer_0[489] ^ layer_0[2001]); 
    assign out[322] = layer_0[1061] ^ layer_0[295]; 
    assign out[323] = layer_0[1313]; 
    assign out[324] = ~(layer_0[587] ^ layer_0[1387]); 
    assign out[325] = ~(layer_0[1847] ^ layer_0[1720]); 
    assign out[326] = layer_0[3318] ^ layer_0[3757]; 
    assign out[327] = ~layer_0[1026] | (layer_0[1026] & layer_0[2945]); 
    assign out[328] = ~layer_0[1963] | (layer_0[1963] & layer_0[547]); 
    assign out[329] = layer_0[3478]; 
    assign out[330] = layer_0[1283] & layer_0[1146]; 
    assign out[331] = layer_0[668] ^ layer_0[3959]; 
    assign out[332] = layer_0[1096] ^ layer_0[2566]; 
    assign out[333] = layer_0[3576] ^ layer_0[993]; 
    assign out[334] = layer_0[1367] ^ layer_0[3127]; 
    assign out[335] = ~(layer_0[2059] ^ layer_0[2281]); 
    assign out[336] = layer_0[442] & ~layer_0[486]; 
    assign out[337] = ~(layer_0[1082] ^ layer_0[239]); 
    assign out[338] = ~(layer_0[1312] | layer_0[3113]); 
    assign out[339] = layer_0[407]; 
    assign out[340] = layer_0[3920] & ~layer_0[2145]; 
    assign out[341] = layer_0[1398] ^ layer_0[2834]; 
    assign out[342] = ~layer_0[1099]; 
    assign out[343] = ~layer_0[954] | (layer_0[1983] & layer_0[954]); 
    assign out[344] = layer_0[127]; 
    assign out[345] = ~layer_0[2967]; 
    assign out[346] = layer_0[2450] ^ layer_0[2431]; 
    assign out[347] = layer_0[423] & ~layer_0[163]; 
    assign out[348] = layer_0[454] ^ layer_0[197]; 
    assign out[349] = layer_0[3257]; 
    assign out[350] = layer_0[1946] ^ layer_0[3693]; 
    assign out[351] = layer_0[1655] & layer_0[2347]; 
    assign out[352] = ~(layer_0[2422] ^ layer_0[2715]); 
    assign out[353] = layer_0[3065] & ~layer_0[693]; 
    assign out[354] = layer_0[1314] & layer_0[1550]; 
    assign out[355] = ~(layer_0[1218] ^ layer_0[3968]); 
    assign out[356] = ~layer_0[2513]; 
    assign out[357] = ~(layer_0[2499] ^ layer_0[1007]); 
    assign out[358] = layer_0[1920] & ~layer_0[3500]; 
    assign out[359] = ~(layer_0[3144] ^ layer_0[309]); 
    assign out[360] = layer_0[662]; 
    assign out[361] = ~(layer_0[2285] ^ layer_0[2401]); 
    assign out[362] = layer_0[1861] ^ layer_0[1119]; 
    assign out[363] = layer_0[1378] ^ layer_0[1245]; 
    assign out[364] = ~layer_0[1358] | (layer_0[818] & layer_0[1358]); 
    assign out[365] = layer_0[1854] ^ layer_0[3908]; 
    assign out[366] = ~(layer_0[2896] ^ layer_0[1560]); 
    assign out[367] = ~(layer_0[966] ^ layer_0[3439]); 
    assign out[368] = ~(layer_0[2387] ^ layer_0[1156]); 
    assign out[369] = layer_0[165]; 
    assign out[370] = ~(layer_0[986] ^ layer_0[822]); 
    assign out[371] = ~layer_0[1104]; 
    assign out[372] = layer_0[1251] ^ layer_0[3613]; 
    assign out[373] = layer_0[3071]; 
    assign out[374] = ~(layer_0[3089] ^ layer_0[1897]); 
    assign out[375] = layer_0[1515] & ~layer_0[1047]; 
    assign out[376] = layer_0[3604] ^ layer_0[177]; 
    assign out[377] = ~(layer_0[3937] ^ layer_0[98]); 
    assign out[378] = layer_0[498] ^ layer_0[3871]; 
    assign out[379] = layer_0[552] & ~layer_0[2226]; 
    assign out[380] = layer_0[3676] & ~layer_0[1181]; 
    assign out[381] = layer_0[402] & ~layer_0[3376]; 
    assign out[382] = layer_0[2256] & ~layer_0[3669]; 
    assign out[383] = ~(layer_0[3410] | layer_0[3928]); 
    assign out[384] = layer_0[2876]; 
    assign out[385] = ~(layer_0[3931] ^ layer_0[753]); 
    assign out[386] = layer_0[1362] ^ layer_0[50]; 
    assign out[387] = layer_0[561] ^ layer_0[2385]; 
    assign out[388] = layer_0[1008] ^ layer_0[2019]; 
    assign out[389] = layer_0[3656] & ~layer_0[3586]; 
    assign out[390] = ~(layer_0[1840] ^ layer_0[3924]); 
    assign out[391] = layer_0[1660] & layer_0[86]; 
    assign out[392] = layer_0[2802]; 
    assign out[393] = layer_0[2612] ^ layer_0[494]; 
    assign out[394] = layer_0[1794] & layer_0[2337]; 
    assign out[395] = ~(layer_0[2375] ^ layer_0[1485]); 
    assign out[396] = layer_0[2887] ^ layer_0[3270]; 
    assign out[397] = layer_0[1422]; 
    assign out[398] = ~(layer_0[1210] | layer_0[1444]); 
    assign out[399] = layer_0[3708] & ~layer_0[618]; 
    assign out[400] = layer_0[1825]; 
    assign out[401] = layer_0[2604]; 
    assign out[402] = ~layer_0[1800]; 
    assign out[403] = ~(layer_0[3388] | layer_0[1851]); 
    assign out[404] = ~(layer_0[1076] ^ layer_0[2306]); 
    assign out[405] = layer_0[2366] & ~layer_0[48]; 
    assign out[406] = layer_0[3519] & ~layer_0[2326]; 
    assign out[407] = layer_0[1091] & ~layer_0[2093]; 
    assign out[408] = layer_0[166]; 
    assign out[409] = ~(layer_0[1589] | layer_0[208]); 
    assign out[410] = ~(layer_0[1406] ^ layer_0[2008]); 
    assign out[411] = ~(layer_0[3508] ^ layer_0[3838]); 
    assign out[412] = ~(layer_0[122] ^ layer_0[1544]); 
    assign out[413] = layer_0[1298] ^ layer_0[199]; 
    assign out[414] = layer_0[1629] ^ layer_0[1178]; 
    assign out[415] = ~(layer_0[3391] | layer_0[2712]); 
    assign out[416] = layer_0[2527] ^ layer_0[2658]; 
    assign out[417] = layer_0[605] & ~layer_0[2294]; 
    assign out[418] = ~layer_0[2685] | (layer_0[2685] & layer_0[3436]); 
    assign out[419] = ~(layer_0[3489] | layer_0[1901]); 
    assign out[420] = layer_0[3936]; 
    assign out[421] = layer_0[2794] & ~layer_0[1914]; 
    assign out[422] = layer_0[2037]; 
    assign out[423] = layer_0[705] & ~layer_0[2307]; 
    assign out[424] = layer_0[1429] & layer_0[404]; 
    assign out[425] = ~(layer_0[3227] | layer_0[1442]); 
    assign out[426] = layer_0[2486]; 
    assign out[427] = layer_0[996]; 
    assign out[428] = layer_0[2361] ^ layer_0[2114]; 
    assign out[429] = ~(layer_0[2423] | layer_0[1950]); 
    assign out[430] = layer_0[2075] & ~layer_0[1235]; 
    assign out[431] = ~layer_0[3662] | (layer_0[3441] & layer_0[3662]); 
    assign out[432] = layer_0[3845] ^ layer_0[592]; 
    assign out[433] = layer_0[1541] & ~layer_0[830]; 
    assign out[434] = layer_0[87] & ~layer_0[1975]; 
    assign out[435] = ~(layer_0[1234] ^ layer_0[271]); 
    assign out[436] = ~layer_0[2550]; 
    assign out[437] = layer_0[2124]; 
    assign out[438] = ~layer_0[2069]; 
    assign out[439] = layer_0[1322] ^ layer_0[679]; 
    assign out[440] = layer_0[1097] ^ layer_0[1495]; 
    assign out[441] = layer_0[1991] & ~layer_0[3430]; 
    assign out[442] = ~(layer_0[3175] & layer_0[2096]); 
    assign out[443] = layer_0[3514] & ~layer_0[2632]; 
    assign out[444] = layer_0[2890] & layer_0[3145]; 
    assign out[445] = ~layer_0[2100]; 
    assign out[446] = layer_0[932] ^ layer_0[385]; 
    assign out[447] = ~(layer_0[126] & layer_0[3372]); 
    assign out[448] = ~(layer_0[109] | layer_0[2525]); 
    assign out[449] = layer_0[389] ^ layer_0[3372]; 
    assign out[450] = layer_0[107] ^ layer_0[1732]; 
    assign out[451] = ~layer_0[1237] | (layer_0[3464] & layer_0[1237]); 
    assign out[452] = layer_0[1324] & ~layer_0[3060]; 
    assign out[453] = layer_0[289] ^ layer_0[292]; 
    assign out[454] = ~(layer_0[642] ^ layer_0[1969]); 
    assign out[455] = layer_0[1794] & layer_0[2510]; 
    assign out[456] = layer_0[3400] ^ layer_0[409]; 
    assign out[457] = layer_0[2933] ^ layer_0[1099]; 
    assign out[458] = ~(layer_0[2275] ^ layer_0[3912]); 
    assign out[459] = layer_0[2116] ^ layer_0[1434]; 
    assign out[460] = layer_0[3992] ^ layer_0[3180]; 
    assign out[461] = layer_0[1344] & layer_0[3872]; 
    assign out[462] = layer_0[957] ^ layer_0[2144]; 
    assign out[463] = layer_0[639]; 
    assign out[464] = layer_0[2944]; 
    assign out[465] = layer_0[2850] ^ layer_0[3795]; 
    assign out[466] = ~layer_0[3948]; 
    assign out[467] = layer_0[3688] & layer_0[1342]; 
    assign out[468] = ~(layer_0[3178] | layer_0[3824]); 
    assign out[469] = layer_0[3981] & layer_0[2252]; 
    assign out[470] = layer_0[236]; 
    assign out[471] = ~layer_0[695]; 
    assign out[472] = layer_0[2387] ^ layer_0[281]; 
    assign out[473] = ~(layer_0[843] | layer_0[763]); 
    assign out[474] = layer_0[3406]; 
    assign out[475] = layer_0[8] & layer_0[2011]; 
    assign out[476] = ~(layer_0[849] | layer_0[692]); 
    assign out[477] = layer_0[1797] ^ layer_0[2817]; 
    assign out[478] = layer_0[1590] & ~layer_0[930]; 
    assign out[479] = layer_0[3097] & ~layer_0[3961]; 
    assign out[480] = ~layer_0[1821]; 
    assign out[481] = layer_0[2163] ^ layer_0[2765]; 
    assign out[482] = ~(layer_0[3149] ^ layer_0[2744]); 
    assign out[483] = layer_0[3046] & layer_0[1376]; 
    assign out[484] = layer_0[570]; 
    assign out[485] = layer_0[3280] & ~layer_0[2717]; 
    assign out[486] = layer_0[1785]; 
    assign out[487] = layer_0[3192] & ~layer_0[1858]; 
    assign out[488] = ~(layer_0[1217] | layer_0[3647]); 
    assign out[489] = ~layer_0[155] | (layer_0[155] & layer_0[1493]); 
    assign out[490] = ~layer_0[581] | (layer_0[581] & layer_0[2086]); 
    assign out[491] = layer_0[2686]; 
    assign out[492] = layer_0[735] & ~layer_0[2709]; 
    assign out[493] = layer_0[3363]; 
    assign out[494] = layer_0[194] ^ layer_0[34]; 
    assign out[495] = layer_0[1805] & ~layer_0[3643]; 
    assign out[496] = layer_0[2458] & ~layer_0[286]; 
    assign out[497] = ~layer_0[2831] | (layer_0[2831] & layer_0[777]); 
    assign out[498] = layer_0[3542] & layer_0[1787]; 
    assign out[499] = layer_0[3177] & ~layer_0[713]; 
    assign out[500] = ~layer_0[1343] | (layer_0[1343] & layer_0[2209]); 
    assign out[501] = layer_0[1143] & ~layer_0[901]; 
    assign out[502] = ~(layer_0[984] ^ layer_0[3610]); 
    assign out[503] = ~(layer_0[3276] ^ layer_0[1539]); 
    assign out[504] = layer_0[368] & ~layer_0[975]; 
    assign out[505] = layer_0[2186] ^ layer_0[1219]; 
    assign out[506] = ~layer_0[1532]; 
    assign out[507] = ~layer_0[3030] | (layer_0[3030] & layer_0[2242]); 
    assign out[508] = layer_0[1925]; 
    assign out[509] = layer_0[865] & ~layer_0[2110]; 
    assign out[510] = ~layer_0[2898]; 
    assign out[511] = ~layer_0[667]; 
    assign out[512] = ~(layer_0[528] ^ layer_0[3599]); 
    assign out[513] = ~layer_0[2515] | (layer_0[2515] & layer_0[3637]); 
    assign out[514] = layer_0[3745] ^ layer_0[3405]; 
    assign out[515] = ~(layer_0[327] ^ layer_0[3001]); 
    assign out[516] = ~(layer_0[3105] ^ layer_0[2438]); 
    assign out[517] = ~(layer_0[929] & layer_0[169]); 
    assign out[518] = ~(layer_0[740] ^ layer_0[654]); 
    assign out[519] = layer_0[1237] & ~layer_0[104]; 
    assign out[520] = layer_0[3887]; 
    assign out[521] = layer_0[1512] ^ layer_0[3277]; 
    assign out[522] = ~(layer_0[340] ^ layer_0[766]); 
    assign out[523] = ~(layer_0[1902] ^ layer_0[2299]); 
    assign out[524] = ~(layer_0[320] & layer_0[3720]); 
    assign out[525] = ~(layer_0[2045] ^ layer_0[1926]); 
    assign out[526] = layer_0[3778] ^ layer_0[1827]; 
    assign out[527] = layer_0[2823] ^ layer_0[3945]; 
    assign out[528] = ~layer_0[3775]; 
    assign out[529] = layer_0[3627] ^ layer_0[1516]; 
    assign out[530] = ~(layer_0[2072] ^ layer_0[14]); 
    assign out[531] = ~layer_0[2487] | (layer_0[2429] & layer_0[2487]); 
    assign out[532] = layer_0[720] ^ layer_0[3763]; 
    assign out[533] = ~(layer_0[2565] ^ layer_0[279]); 
    assign out[534] = ~layer_0[795] | (layer_0[795] & layer_0[1310]); 
    assign out[535] = ~(layer_0[1535] ^ layer_0[76]); 
    assign out[536] = ~layer_0[2737]; 
    assign out[537] = layer_0[3773]; 
    assign out[538] = ~layer_0[1003]; 
    assign out[539] = layer_0[2295] ^ layer_0[1753]; 
    assign out[540] = layer_0[59] ^ layer_0[3077]; 
    assign out[541] = ~(layer_0[471] ^ layer_0[2042]); 
    assign out[542] = ~layer_0[784]; 
    assign out[543] = layer_0[2596] ^ layer_0[1832]; 
    assign out[544] = ~(layer_0[3240] ^ layer_0[1741]); 
    assign out[545] = layer_0[3039] ^ layer_0[234]; 
    assign out[546] = ~layer_0[2815]; 
    assign out[547] = ~layer_0[3244]; 
    assign out[548] = layer_0[890] | layer_0[1414]; 
    assign out[549] = ~layer_0[282]; 
    assign out[550] = ~layer_0[3359]; 
    assign out[551] = ~(layer_0[1154] ^ layer_0[1731]); 
    assign out[552] = ~layer_0[142]; 
    assign out[553] = layer_0[3428] & ~layer_0[460]; 
    assign out[554] = ~(layer_0[3891] & layer_0[2980]); 
    assign out[555] = layer_0[780] ^ layer_0[1119]; 
    assign out[556] = layer_0[2993]; 
    assign out[557] = ~(layer_0[3825] ^ layer_0[1098]); 
    assign out[558] = layer_0[3271] ^ layer_0[3735]; 
    assign out[559] = layer_0[2670]; 
    assign out[560] = ~layer_0[3759]; 
    assign out[561] = ~(layer_0[1457] & layer_0[315]); 
    assign out[562] = ~(layer_0[579] ^ layer_0[3964]); 
    assign out[563] = ~layer_0[3263]; 
    assign out[564] = ~layer_0[1169] | (layer_0[1169] & layer_0[564]); 
    assign out[565] = layer_0[3902] ^ layer_0[1]; 
    assign out[566] = layer_0[2311] ^ layer_0[23]; 
    assign out[567] = layer_0[1172] | layer_0[1443]; 
    assign out[568] = layer_0[2324] & layer_0[3343]; 
    assign out[569] = ~(layer_0[3650] ^ layer_0[3184]); 
    assign out[570] = layer_0[3619] & ~layer_0[1713]; 
    assign out[571] = ~(layer_0[3962] ^ layer_0[655]); 
    assign out[572] = ~(layer_0[1221] ^ layer_0[1381]); 
    assign out[573] = ~(layer_0[2339] & layer_0[2958]); 
    assign out[574] = layer_0[2215] ^ layer_0[1075]; 
    assign out[575] = layer_0[2204] ^ layer_0[3915]; 
    assign out[576] = layer_0[2493] | layer_0[1781]; 
    assign out[577] = layer_0[1880] ^ layer_0[2736]; 
    assign out[578] = ~layer_0[517]; 
    assign out[579] = ~(layer_0[1078] ^ layer_0[2118]); 
    assign out[580] = layer_0[2542] ^ layer_0[369]; 
    assign out[581] = ~(layer_0[941] ^ layer_0[3098]); 
    assign out[582] = layer_0[3471] ^ layer_0[1819]; 
    assign out[583] = layer_0[3436]; 
    assign out[584] = layer_0[2205]; 
    assign out[585] = layer_0[2120] ^ layer_0[1980]; 
    assign out[586] = ~(layer_0[1917] ^ layer_0[962]); 
    assign out[587] = layer_0[11] ^ layer_0[829]; 
    assign out[588] = layer_0[3534] ^ layer_0[261]; 
    assign out[589] = ~(layer_0[1117] & layer_0[2895]); 
    assign out[590] = layer_0[3984] ^ layer_0[1265]; 
    assign out[591] = ~layer_0[3893]; 
    assign out[592] = ~(layer_0[2767] ^ layer_0[2820]); 
    assign out[593] = layer_0[1106] ^ layer_0[3518]; 
    assign out[594] = layer_0[3148] & ~layer_0[3649]; 
    assign out[595] = layer_0[2804] ^ layer_0[3877]; 
    assign out[596] = layer_0[1465] ^ layer_0[3917]; 
    assign out[597] = layer_0[3052] ^ layer_0[532]; 
    assign out[598] = ~layer_0[2553] | (layer_0[2553] & layer_0[3886]); 
    assign out[599] = layer_0[738] ^ layer_0[3726]; 
    assign out[600] = ~(layer_0[2605] ^ layer_0[767]); 
    assign out[601] = layer_0[216] & ~layer_0[1867]; 
    assign out[602] = ~(layer_0[1273] ^ layer_0[3229]); 
    assign out[603] = ~(layer_0[2078] ^ layer_0[3607]); 
    assign out[604] = ~(layer_0[1250] ^ layer_0[1124]); 
    assign out[605] = layer_0[158] ^ layer_0[3851]; 
    assign out[606] = ~(layer_0[3986] & layer_0[1070]); 
    assign out[607] = layer_0[1531]; 
    assign out[608] = ~layer_0[1823] | (layer_0[1095] & layer_0[1823]); 
    assign out[609] = ~(layer_0[1519] ^ layer_0[3316]); 
    assign out[610] = ~layer_0[2305]; 
    assign out[611] = layer_0[2213]; 
    assign out[612] = layer_0[1450] ^ layer_0[2111]; 
    assign out[613] = ~(layer_0[814] | layer_0[1190]); 
    assign out[614] = layer_0[2883] ^ layer_0[3950]; 
    assign out[615] = ~(layer_0[2496] ^ layer_0[3063]); 
    assign out[616] = layer_0[836] ^ layer_0[80]; 
    assign out[617] = layer_0[2552] & ~layer_0[2483]; 
    assign out[618] = layer_0[1376] ^ layer_0[3176]; 
    assign out[619] = layer_0[3512] ^ layer_0[1205]; 
    assign out[620] = layer_0[3570] ^ layer_0[2755]; 
    assign out[621] = layer_0[1739] & ~layer_0[2666]; 
    assign out[622] = layer_0[2910] | layer_0[2377]; 
    assign out[623] = ~layer_0[3503]; 
    assign out[624] = layer_0[1056]; 
    assign out[625] = ~layer_0[3409] | (layer_0[3109] & layer_0[3409]); 
    assign out[626] = layer_0[935]; 
    assign out[627] = layer_0[625] | layer_0[1987]; 
    assign out[628] = ~layer_0[3029]; 
    assign out[629] = layer_0[3224] ^ layer_0[3141]; 
    assign out[630] = layer_0[3797] | layer_0[1651]; 
    assign out[631] = ~(layer_0[2086] ^ layer_0[1348]); 
    assign out[632] = layer_0[2653] & ~layer_0[3841]; 
    assign out[633] = layer_0[2427] ^ layer_0[230]; 
    assign out[634] = layer_0[3833]; 
    assign out[635] = ~(layer_0[684] ^ layer_0[3587]); 
    assign out[636] = ~(layer_0[1596] ^ layer_0[1050]); 
    assign out[637] = layer_0[3490]; 
    assign out[638] = layer_0[1790] ^ layer_0[638]; 
    assign out[639] = layer_0[2459] ^ layer_0[2091]; 
    assign out[640] = layer_0[1752] ^ layer_0[747]; 
    assign out[641] = layer_0[1866]; 
    assign out[642] = ~layer_0[1727] | (layer_0[1200] & layer_0[1727]); 
    assign out[643] = ~layer_0[303]; 
    assign out[644] = layer_0[1554] | layer_0[2320]; 
    assign out[645] = ~layer_0[3578]; 
    assign out[646] = ~layer_0[1656]; 
    assign out[647] = ~(layer_0[2280] & layer_0[2470]); 
    assign out[648] = ~(layer_0[2468] ^ layer_0[1033]); 
    assign out[649] = layer_0[257] & ~layer_0[3217]; 
    assign out[650] = layer_0[2873] ^ layer_0[1157]; 
    assign out[651] = layer_0[2733]; 
    assign out[652] = layer_0[2500] | layer_0[190]; 
    assign out[653] = ~(layer_0[1] ^ layer_0[907]); 
    assign out[654] = ~layer_0[3635]; 
    assign out[655] = ~(layer_0[105] & layer_0[104]); 
    assign out[656] = layer_0[3772] & layer_0[3093]; 
    assign out[657] = ~(layer_0[1867] & layer_0[3156]); 
    assign out[658] = ~layer_0[3243] | (layer_0[3243] & layer_0[680]); 
    assign out[659] = ~(layer_0[2860] ^ layer_0[1316]); 
    assign out[660] = layer_0[1384] ^ layer_0[454]; 
    assign out[661] = ~layer_0[2538]; 
    assign out[662] = ~layer_0[1698]; 
    assign out[663] = ~layer_0[821]; 
    assign out[664] = layer_0[2738] ^ layer_0[85]; 
    assign out[665] = ~(layer_0[1862] ^ layer_0[1567]); 
    assign out[666] = ~layer_0[361]; 
    assign out[667] = layer_0[3138] & ~layer_0[3629]; 
    assign out[668] = ~layer_0[3502]; 
    assign out[669] = ~(layer_0[1723] & layer_0[1609]); 
    assign out[670] = ~(layer_0[3542] ^ layer_0[1918]); 
    assign out[671] = layer_0[2553] ^ layer_0[2125]; 
    assign out[672] = layer_0[3679] ^ layer_0[2260]; 
    assign out[673] = layer_0[1240]; 
    assign out[674] = ~layer_0[953]; 
    assign out[675] = layer_0[1696] ^ layer_0[589]; 
    assign out[676] = ~(layer_0[980] ^ layer_0[1829]); 
    assign out[677] = layer_0[2927] & ~layer_0[415]; 
    assign out[678] = layer_0[2507] & ~layer_0[60]; 
    assign out[679] = ~layer_0[3461]; 
    assign out[680] = layer_0[2059]; 
    assign out[681] = layer_0[1302]; 
    assign out[682] = ~(layer_0[2789] ^ layer_0[2087]); 
    assign out[683] = layer_0[3417] ^ layer_0[2905]; 
    assign out[684] = ~(layer_0[77] ^ layer_0[968]); 
    assign out[685] = ~layer_0[787]; 
    assign out[686] = layer_0[3116] ^ layer_0[159]; 
    assign out[687] = layer_0[1403] ^ layer_0[2783]; 
    assign out[688] = ~layer_0[1081]; 
    assign out[689] = layer_0[3183]; 
    assign out[690] = ~(layer_0[231] ^ layer_0[2900]); 
    assign out[691] = ~(layer_0[1490] ^ layer_0[748]); 
    assign out[692] = layer_0[2589]; 
    assign out[693] = layer_0[1968] ^ layer_0[3612]; 
    assign out[694] = ~(layer_0[2258] & layer_0[998]); 
    assign out[695] = ~layer_0[3310] | (layer_0[19] & layer_0[3310]); 
    assign out[696] = ~(layer_0[896] | layer_0[3347]); 
    assign out[697] = ~(layer_0[1029] ^ layer_0[1954]); 
    assign out[698] = ~(layer_0[3278] ^ layer_0[2497]); 
    assign out[699] = ~(layer_0[772] ^ layer_0[2514]); 
    assign out[700] = layer_0[1762] ^ layer_0[1917]; 
    assign out[701] = layer_0[2302] ^ layer_0[2536]; 
    assign out[702] = layer_0[858] ^ layer_0[2556]; 
    assign out[703] = ~layer_0[228] | (layer_0[2191] & layer_0[228]); 
    assign out[704] = layer_0[3284] & ~layer_0[1581]; 
    assign out[705] = ~(layer_0[2682] & layer_0[3407]); 
    assign out[706] = layer_0[870] & layer_0[2002]; 
    assign out[707] = layer_0[3524] ^ layer_0[2849]; 
    assign out[708] = ~(layer_0[2363] ^ layer_0[3266]); 
    assign out[709] = layer_0[1173] & ~layer_0[686]; 
    assign out[710] = layer_0[1838]; 
    assign out[711] = layer_0[3314]; 
    assign out[712] = ~(layer_0[2864] ^ layer_0[3380]); 
    assign out[713] = layer_0[1527] ^ layer_0[2444]; 
    assign out[714] = ~layer_0[3090]; 
    assign out[715] = ~(layer_0[3785] ^ layer_0[586]); 
    assign out[716] = ~(layer_0[3294] & layer_0[1640]); 
    assign out[717] = layer_0[895] & layer_0[3167]; 
    assign out[718] = ~(layer_0[1778] ^ layer_0[3561]); 
    assign out[719] = layer_0[3521] & ~layer_0[3540]; 
    assign out[720] = ~(layer_0[509] ^ layer_0[621]); 
    assign out[721] = ~(layer_0[3402] ^ layer_0[3969]); 
    assign out[722] = layer_0[3768]; 
    assign out[723] = layer_0[3070] | layer_0[3120]; 
    assign out[724] = ~(layer_0[3786] ^ layer_0[367]); 
    assign out[725] = layer_0[874] & ~layer_0[1463]; 
    assign out[726] = ~(layer_0[2649] ^ layer_0[1915]); 
    assign out[727] = ~layer_0[2615] | (layer_0[2615] & layer_0[235]); 
    assign out[728] = layer_0[1427]; 
    assign out[729] = layer_0[1504] | layer_0[2975]; 
    assign out[730] = ~(layer_0[401] & layer_0[2719]); 
    assign out[731] = layer_0[2751] ^ layer_0[2786]; 
    assign out[732] = layer_0[1970] & ~layer_0[3680]; 
    assign out[733] = ~(layer_0[1184] | layer_0[53]); 
    assign out[734] = layer_0[1699] & ~layer_0[2750]; 
    assign out[735] = layer_0[3932] ^ layer_0[3397]; 
    assign out[736] = layer_0[46] ^ layer_0[287]; 
    assign out[737] = layer_0[2598]; 
    assign out[738] = ~(layer_0[2623] ^ layer_0[978]); 
    assign out[739] = ~layer_0[2102] | (layer_0[2102] & layer_0[3101]); 
    assign out[740] = ~(layer_0[2758] & layer_0[193]); 
    assign out[741] = ~layer_0[2530]; 
    assign out[742] = ~(layer_0[711] ^ layer_0[1182]); 
    assign out[743] = ~(layer_0[558] ^ layer_0[1909]); 
    assign out[744] = ~(layer_0[3468] ^ layer_0[1373]); 
    assign out[745] = ~layer_0[1700]; 
    assign out[746] = layer_0[1688] & ~layer_0[2161]; 
    assign out[747] = ~layer_0[3844]; 
    assign out[748] = ~(layer_0[1999] ^ layer_0[2964]); 
    assign out[749] = layer_0[1042] & ~layer_0[2222]; 
    assign out[750] = ~(layer_0[3522] ^ layer_0[1127]); 
    assign out[751] = layer_0[1831]; 
    assign out[752] = layer_0[539] & layer_0[1734]; 
    assign out[753] = layer_0[2561] & layer_0[2498]; 
    assign out[754] = layer_0[2701] ^ layer_0[992]; 
    assign out[755] = ~layer_0[2199] | (layer_0[191] & layer_0[2199]); 
    assign out[756] = ~(layer_0[2979] ^ layer_0[242]); 
    assign out[757] = ~layer_0[1339]; 
    assign out[758] = layer_0[733] ^ layer_0[1228]; 
    assign out[759] = ~layer_0[1132]; 
    assign out[760] = layer_0[3717]; 
    assign out[761] = ~layer_0[881] | (layer_0[2412] & layer_0[881]); 
    assign out[762] = ~layer_0[1760] | (layer_0[2662] & layer_0[1760]); 
    assign out[763] = ~layer_0[1646] | (layer_0[1646] & layer_0[2068]); 
    assign out[764] = layer_0[3099] ^ layer_0[2690]; 
    assign out[765] = ~layer_0[2576]; 
    assign out[766] = layer_0[3904] ^ layer_0[2064]; 
    assign out[767] = layer_0[2126]; 
    assign out[768] = layer_0[2082]; 
    assign out[769] = ~(layer_0[827] & layer_0[222]); 
    assign out[770] = layer_0[2885] & ~layer_0[2032]; 
    assign out[771] = ~(layer_0[3361] ^ layer_0[943]); 
    assign out[772] = ~layer_0[54] | (layer_0[1439] & layer_0[54]); 
    assign out[773] = ~layer_0[2982] | (layer_0[2982] & layer_0[3481]); 
    assign out[774] = ~(layer_0[1478] | layer_0[2939]); 
    assign out[775] = ~layer_0[641] | (layer_0[2752] & layer_0[641]); 
    assign out[776] = ~layer_0[3198]; 
    assign out[777] = ~(layer_0[2330] & layer_0[956]); 
    assign out[778] = layer_0[2654] ^ layer_0[1967]; 
    assign out[779] = layer_0[1649] & ~layer_0[357]; 
    assign out[780] = ~layer_0[1671] | (layer_0[3925] & layer_0[1671]); 
    assign out[781] = layer_0[333] & ~layer_0[572]; 
    assign out[782] = layer_0[1631] & layer_0[683]; 
    assign out[783] = layer_0[1514] ^ layer_0[2047]; 
    assign out[784] = layer_0[908] & ~layer_0[3338]; 
    assign out[785] = ~(layer_0[2652] | layer_0[2325]); 
    assign out[786] = ~(layer_0[1176] ^ layer_0[1716]); 
    assign out[787] = ~layer_0[568] | (layer_0[3365] & layer_0[568]); 
    assign out[788] = layer_0[3429] ^ layer_0[732]; 
    assign out[789] = layer_0[701] ^ layer_0[1114]; 
    assign out[790] = ~(layer_0[2529] ^ layer_0[1263]); 
    assign out[791] = layer_0[1932] & ~layer_0[565]; 
    assign out[792] = ~(layer_0[2317] ^ layer_0[66]); 
    assign out[793] = ~layer_0[559] | (layer_0[1835] & layer_0[559]); 
    assign out[794] = layer_0[384] & layer_0[1462]; 
    assign out[795] = layer_0[3783] ^ layer_0[3237]; 
    assign out[796] = ~(layer_0[937] & layer_0[3182]); 
    assign out[797] = ~layer_0[827] | (layer_0[2655] & layer_0[827]); 
    assign out[798] = layer_0[285] & ~layer_0[3271]; 
    assign out[799] = layer_0[108]; 
    assign out[800] = ~layer_0[1349]; 
    assign out[801] = ~(layer_0[1815] ^ layer_0[3130]); 
    assign out[802] = layer_0[3718] & ~layer_0[2039]; 
    assign out[803] = ~(layer_0[2491] ^ layer_0[205]); 
    assign out[804] = layer_0[2211] ^ layer_0[3907]; 
    assign out[805] = layer_0[1789] & layer_0[1605]; 
    assign out[806] = ~(layer_0[3039] | layer_0[338]); 
    assign out[807] = ~(layer_0[1038] ^ layer_0[1385]); 
    assign out[808] = layer_0[166]; 
    assign out[809] = ~(layer_0[2687] ^ layer_0[32]); 
    assign out[810] = layer_0[3335] ^ layer_0[3517]; 
    assign out[811] = layer_0[1304] ^ layer_0[2356]; 
    assign out[812] = ~layer_0[1148] | (layer_0[1148] & layer_0[3933]); 
    assign out[813] = ~(layer_0[3967] ^ layer_0[3741]); 
    assign out[814] = layer_0[3412] & layer_0[2511]; 
    assign out[815] = ~(layer_0[1736] ^ layer_0[21]); 
    assign out[816] = layer_0[322] | layer_0[2073]; 
    assign out[817] = layer_0[2766] ^ layer_0[2101]; 
    assign out[818] = layer_0[2370]; 
    assign out[819] = ~layer_0[563]; 
    assign out[820] = layer_0[2003] & layer_0[1041]; 
    assign out[821] = ~layer_0[3085]; 
    assign out[822] = ~layer_0[602]; 
    assign out[823] = layer_0[2551] & layer_0[3514]; 
    assign out[824] = ~(layer_0[1601] ^ layer_0[875]); 
    assign out[825] = ~(layer_0[3704] ^ layer_0[1141]); 
    assign out[826] = ~layer_0[2254]; 
    assign out[827] = layer_0[2348] & ~layer_0[3636]; 
    assign out[828] = layer_0[2960] | layer_0[1962]; 
    assign out[829] = layer_0[2121] ^ layer_0[1799]; 
    assign out[830] = ~layer_0[3993]; 
    assign out[831] = ~(layer_0[999] ^ layer_0[2277]); 
    assign out[832] = ~(layer_0[3557] ^ layer_0[2841]); 
    assign out[833] = layer_0[1167] ^ layer_0[2561]; 
    assign out[834] = layer_0[1563] & ~layer_0[1935]; 
    assign out[835] = layer_0[230] & ~layer_0[2855]; 
    assign out[836] = ~(layer_0[1275] ^ layer_0[2180]); 
    assign out[837] = layer_0[809] ^ layer_0[774]; 
    assign out[838] = ~(layer_0[135] ^ layer_0[2673]); 
    assign out[839] = ~layer_0[81]; 
    assign out[840] = layer_0[3589]; 
    assign out[841] = layer_0[426] ^ layer_0[1126]; 
    assign out[842] = layer_0[853] ^ layer_0[3336]; 
    assign out[843] = ~layer_0[1006]; 
    assign out[844] = layer_0[2122] & ~layer_0[420]; 
    assign out[845] = layer_0[1460] ^ layer_0[1884]; 
    assign out[846] = layer_0[2092]; 
    assign out[847] = ~layer_0[1071] | (layer_0[1071] & layer_0[2288]); 
    assign out[848] = ~layer_0[253] | (layer_0[354] & layer_0[253]); 
    assign out[849] = ~(layer_0[3940] ^ layer_0[3325]); 
    assign out[850] = ~layer_0[3861]; 
    assign out[851] = layer_0[2951] & ~layer_0[3443]; 
    assign out[852] = layer_0[2191] & ~layer_0[9]; 
    assign out[853] = layer_0[3139] ^ layer_0[1480]; 
    assign out[854] = ~layer_0[2032] | (layer_0[1984] & layer_0[2032]); 
    assign out[855] = layer_0[347] ^ layer_0[1530]; 
    assign out[856] = layer_0[1885]; 
    assign out[857] = ~layer_0[3018] | (layer_0[3018] & layer_0[2889]); 
    assign out[858] = layer_0[27] ^ layer_0[3106]; 
    assign out[859] = layer_0[2357] & ~layer_0[1285]; 
    assign out[860] = layer_0[2636]; 
    assign out[861] = ~layer_0[3181]; 
    assign out[862] = ~(layer_0[33] ^ layer_0[3746]); 
    assign out[863] = layer_0[2697] & layer_0[2446]; 
    assign out[864] = layer_0[192] ^ layer_0[1012]; 
    assign out[865] = layer_0[3579] & ~layer_0[149]; 
    assign out[866] = ~(layer_0[1397] ^ layer_0[77]); 
    assign out[867] = ~(layer_0[1374] ^ layer_0[3603]); 
    assign out[868] = ~(layer_0[2652] ^ layer_0[1092]); 
    assign out[869] = ~layer_0[825] | (layer_0[925] & layer_0[825]); 
    assign out[870] = ~(layer_0[739] ^ layer_0[2300]); 
    assign out[871] = layer_0[125] | layer_0[782]; 
    assign out[872] = layer_0[2136] & layer_0[3885]; 
    assign out[873] = ~layer_0[841]; 
    assign out[874] = layer_0[3536] ^ layer_0[2160]; 
    assign out[875] = ~(layer_0[1177] ^ layer_0[2537]); 
    assign out[876] = layer_0[2599]; 
    assign out[877] = layer_0[1346] | layer_0[816]; 
    assign out[878] = ~layer_0[1123] | (layer_0[1123] & layer_0[2801]); 
    assign out[879] = layer_0[1515] & ~layer_0[1269]; 
    assign out[880] = layer_0[3577] ^ layer_0[1642]; 
    assign out[881] = layer_0[838]; 
    assign out[882] = ~(layer_0[2506] & layer_0[2539]); 
    assign out[883] = ~layer_0[656]; 
    assign out[884] = layer_0[3994] & ~layer_0[671]; 
    assign out[885] = layer_0[3503] & ~layer_0[3325]; 
    assign out[886] = ~layer_0[3480]; 
    assign out[887] = layer_0[1795] & ~layer_0[1553]; 
    assign out[888] = layer_0[1947] & layer_0[3784]; 
    assign out[889] = layer_0[299] ^ layer_0[3256]; 
    assign out[890] = ~(layer_0[1042] & layer_0[1152]); 
    assign out[891] = ~layer_0[689]; 
    assign out[892] = layer_0[2373] ^ layer_0[677]; 
    assign out[893] = layer_0[2725]; 
    assign out[894] = ~layer_0[624] | (layer_0[624] & layer_0[726]); 
    assign out[895] = layer_0[581] ^ layer_0[3721]; 
    assign out[896] = ~(layer_0[773] | layer_0[2619]); 
    assign out[897] = ~(layer_0[2842] | layer_0[48]); 
    assign out[898] = ~(layer_0[2164] ^ layer_0[3790]); 
    assign out[899] = ~layer_0[3374] | (layer_0[1422] & layer_0[3374]); 
    assign out[900] = ~layer_0[3911] | (layer_0[2372] & layer_0[3911]); 
    assign out[901] = layer_0[1325] ^ layer_0[1764]; 
    assign out[902] = layer_0[2728]; 
    assign out[903] = layer_0[1330] | layer_0[1657]; 
    assign out[904] = layer_0[3664] ^ layer_0[2935]; 
    assign out[905] = layer_0[3107]; 
    assign out[906] = ~(layer_0[2577] ^ layer_0[1538]); 
    assign out[907] = layer_0[2567]; 
    assign out[908] = layer_0[1786] & layer_0[2511]; 
    assign out[909] = ~(layer_0[427] ^ layer_0[2665]); 
    assign out[910] = ~(layer_0[3979] & layer_0[892]); 
    assign out[911] = ~layer_0[3592] | (layer_0[3839] & layer_0[3592]); 
    assign out[912] = ~layer_0[3600] | (layer_0[105] & layer_0[3600]); 
    assign out[913] = ~layer_0[831]; 
    assign out[914] = layer_0[3487] & ~layer_0[3223]; 
    assign out[915] = ~layer_0[2754] | (layer_0[2754] & layer_0[2479]); 
    assign out[916] = ~(layer_0[1199] ^ layer_0[2268]); 
    assign out[917] = ~(layer_0[2253] ^ layer_0[2718]); 
    assign out[918] = ~layer_0[2770] | (layer_0[2984] & layer_0[2770]); 
    assign out[919] = layer_0[1619] ^ layer_0[2416]; 
    assign out[920] = layer_0[1658] & ~layer_0[3056]; 
    assign out[921] = layer_0[3719] ^ layer_0[489]; 
    assign out[922] = ~layer_0[1933] | (layer_0[1933] & layer_0[2658]); 
    assign out[923] = ~(layer_0[2790] ^ layer_0[2697]); 
    assign out[924] = layer_0[1412] & ~layer_0[3787]; 
    assign out[925] = ~(layer_0[210] | layer_0[572]); 
    assign out[926] = layer_0[3426] ^ layer_0[3049]; 
    assign out[927] = layer_0[1886]; 
    assign out[928] = ~(layer_0[1332] ^ layer_0[2680]); 
    assign out[929] = layer_0[793] ^ layer_0[1994]; 
    assign out[930] = ~(layer_0[3665] ^ layer_0[1458]); 
    assign out[931] = ~(layer_0[2296] ^ layer_0[3632]); 
    assign out[932] = layer_0[2405] & layer_0[2994]; 
    assign out[933] = ~(layer_0[1930] ^ layer_0[2795]); 
    assign out[934] = ~layer_0[646]; 
    assign out[935] = layer_0[3868] ^ layer_0[859]; 
    assign out[936] = layer_0[3586] ^ layer_0[3906]; 
    assign out[937] = layer_0[1528]; 
    assign out[938] = layer_0[1937] & ~layer_0[3387]; 
    assign out[939] = layer_0[512] & ~layer_0[1611]; 
    assign out[940] = layer_0[526] ^ layer_0[1600]; 
    assign out[941] = ~(layer_0[1220] ^ layer_0[2839]); 
    assign out[942] = ~(layer_0[493] ^ layer_0[2175]); 
    assign out[943] = layer_0[3590] & layer_0[1937]; 
    assign out[944] = layer_0[2415] & layer_0[436]; 
    assign out[945] = layer_0[3843] & layer_0[1052]; 
    assign out[946] = ~layer_0[3260] | (layer_0[1014] & layer_0[3260]); 
    assign out[947] = ~(layer_0[1725] ^ layer_0[2557]); 
    assign out[948] = ~layer_0[1145]; 
    assign out[949] = layer_0[696] & ~layer_0[1714]; 
    assign out[950] = ~layer_0[1636]; 
    assign out[951] = layer_0[3233] & layer_0[1682]; 
    assign out[952] = layer_0[2237]; 
    assign out[953] = layer_0[3509]; 
    assign out[954] = ~(layer_0[274] | layer_0[595]); 
    assign out[955] = layer_0[511] ^ layer_0[3566]; 
    assign out[956] = layer_0[3568] & ~layer_0[2140]; 
    assign out[957] = layer_0[1907] & ~layer_0[3299]; 
    assign out[958] = ~(layer_0[1093] | layer_0[3852]); 
    assign out[959] = ~layer_0[140]; 
    assign out[960] = ~(layer_0[3771] | layer_0[3540]); 
    assign out[961] = layer_0[3122] & layer_0[3467]; 
    assign out[962] = ~layer_0[338]; 
    assign out[963] = layer_0[3595] ^ layer_0[1116]; 
    assign out[964] = ~layer_0[2865]; 
    assign out[965] = ~layer_0[1248] | (layer_0[1248] & layer_0[504]); 
    assign out[966] = layer_0[1236] & ~layer_0[2282]; 
    assign out[967] = ~(layer_0[1309] ^ layer_0[2098]); 
    assign out[968] = ~(layer_0[3322] | layer_0[3789]); 
    assign out[969] = layer_0[850] & layer_0[3168]; 
    assign out[970] = layer_0[870]; 
    assign out[971] = layer_0[3283] | layer_0[919]; 
    assign out[972] = ~(layer_0[3320] ^ layer_0[2112]); 
    assign out[973] = ~(layer_0[403] ^ layer_0[2916]); 
    assign out[974] = ~(layer_0[3624] | layer_0[1285]); 
    assign out[975] = layer_0[356] ^ layer_0[364]; 
    assign out[976] = ~(layer_0[3147] ^ layer_0[267]); 
    assign out[977] = layer_0[2718] ^ layer_0[2172]; 
    assign out[978] = ~(layer_0[355] ^ layer_0[1347]); 
    assign out[979] = ~(layer_0[2522] ^ layer_0[1461]); 
    assign out[980] = ~(layer_0[2974] ^ layer_0[1801]); 
    assign out[981] = ~layer_0[3064] | (layer_0[3812] & layer_0[3064]); 
    assign out[982] = ~(layer_0[3595] ^ layer_0[1868]); 
    assign out[983] = layer_0[527] | layer_0[3689]; 
    assign out[984] = layer_0[3488] & ~layer_0[3624]; 
    assign out[985] = layer_0[3125] ^ layer_0[2273]; 
    assign out[986] = ~(layer_0[3707] ^ layer_0[1451]); 
    assign out[987] = layer_0[3096] ^ layer_0[562]; 
    assign out[988] = ~layer_0[3955]; 
    assign out[989] = ~(layer_0[3618] ^ layer_0[2562]); 
    assign out[990] = layer_0[3760] ^ layer_0[2559]; 
    assign out[991] = ~layer_0[1135] | (layer_0[1135] & layer_0[967]); 
    assign out[992] = ~(layer_0[3922] ^ layer_0[1483]); 
    assign out[993] = ~(layer_0[2844] ^ layer_0[3368]); 
    assign out[994] = ~(layer_0[3118] ^ layer_0[1583]); 
    assign out[995] = ~layer_0[2018] | (layer_0[1390] & layer_0[2018]); 
    assign out[996] = layer_0[1686] | layer_0[3544]; 
    assign out[997] = layer_0[1506] & ~layer_0[3699]; 
    assign out[998] = ~layer_0[1887]; 
    assign out[999] = ~(layer_0[3538] | layer_0[1365]); 
    assign out[1000] = ~layer_0[3255] | (layer_0[1281] & layer_0[3255]); 
    assign out[1001] = layer_0[1711] ^ layer_0[2477]; 
    assign out[1002] = ~layer_0[210]; 
    assign out[1003] = layer_0[2526] ^ layer_0[1961]; 
    assign out[1004] = ~(layer_0[444] ^ layer_0[3193]); 
    assign out[1005] = ~(layer_0[2990] ^ layer_0[3408]); 
    assign out[1006] = ~(layer_0[258] ^ layer_0[2618]); 
    assign out[1007] = layer_0[1044] ^ layer_0[3946]; 
    assign out[1008] = ~(layer_0[3304] ^ layer_0[3914]); 
    assign out[1009] = ~(layer_0[609] ^ layer_0[2297]); 
    assign out[1010] = layer_0[144] ^ layer_0[1945]; 
    assign out[1011] = ~(layer_0[392] ^ layer_0[3164]); 
    assign out[1012] = ~(layer_0[3505] ^ layer_0[1751]); 
    assign out[1013] = layer_0[3380] ^ layer_0[2223]; 
    assign out[1014] = layer_0[2051] ^ layer_0[3914]; 
    assign out[1015] = layer_0[815] ^ layer_0[360]; 
    assign out[1016] = layer_0[1922] | layer_0[416]; 
    assign out[1017] = ~(layer_0[2168] ^ layer_0[906]); 
    assign out[1018] = layer_0[3983]; 
    assign out[1019] = layer_0[2149] ^ layer_0[3432]; 
    assign out[1020] = layer_0[418]; 
    assign out[1021] = ~layer_0[1591] | (layer_0[1591] & layer_0[3901]); 
    assign out[1022] = ~(layer_0[2880] ^ layer_0[677]); 
    assign out[1023] = layer_0[2827]; 
    assign out[1024] = layer_0[651] ^ layer_0[3776]; 
    assign out[1025] = ~(layer_0[1197] ^ layer_0[1460]); 
    assign out[1026] = layer_0[1141] & ~layer_0[3267]; 
    assign out[1027] = layer_0[1718] ^ layer_0[3840]; 
    assign out[1028] = layer_0[200] ^ layer_0[1202]; 
    assign out[1029] = layer_0[1764]; 
    assign out[1030] = layer_0[1521] & layer_0[3169]; 
    assign out[1031] = ~layer_0[3711] | (layer_0[409] & layer_0[3711]); 
    assign out[1032] = layer_0[2184] & ~layer_0[1733]; 
    assign out[1033] = layer_0[2535] & layer_0[2268]; 
    assign out[1034] = layer_0[1367]; 
    assign out[1035] = ~layer_0[2378]; 
    assign out[1036] = ~layer_0[3645]; 
    assign out[1037] = ~(layer_0[91] ^ layer_0[2921]); 
    assign out[1038] = ~layer_0[476]; 
    assign out[1039] = ~layer_0[1352] | (layer_0[691] & layer_0[1352]); 
    assign out[1040] = layer_0[1194] ^ layer_0[2972]; 
    assign out[1041] = ~layer_0[1361]; 
    assign out[1042] = layer_0[2859]; 
    assign out[1043] = layer_0[1694]; 
    assign out[1044] = ~layer_0[1547] | (layer_0[1473] & layer_0[1547]); 
    assign out[1045] = ~layer_0[1782]; 
    assign out[1046] = layer_0[1008] & ~layer_0[2795]; 
    assign out[1047] = ~(layer_0[3425] ^ layer_0[276]); 
    assign out[1048] = ~(layer_0[2840] ^ layer_0[178]); 
    assign out[1049] = ~(layer_0[1067] ^ layer_0[1157]); 
    assign out[1050] = ~layer_0[2166]; 
    assign out[1051] = ~(layer_0[1498] & layer_0[45]); 
    assign out[1052] = layer_0[1428] | layer_0[202]; 
    assign out[1053] = layer_0[297] ^ layer_0[52]; 
    assign out[1054] = layer_0[2094] | layer_0[1744]; 
    assign out[1055] = ~layer_0[3467]; 
    assign out[1056] = layer_0[2913] ^ layer_0[1616]; 
    assign out[1057] = ~layer_0[2066]; 
    assign out[1058] = ~(layer_0[3151] ^ layer_0[3672]); 
    assign out[1059] = ~(layer_0[2110] ^ layer_0[1352]); 
    assign out[1060] = layer_0[3856] ^ layer_0[965]; 
    assign out[1061] = ~layer_0[3906] | (layer_0[3906] & layer_0[2151]); 
    assign out[1062] = ~(layer_0[3342] & layer_0[3073]); 
    assign out[1063] = ~(layer_0[542] ^ layer_0[416]); 
    assign out[1064] = ~(layer_0[2448] ^ layer_0[802]); 
    assign out[1065] = ~(layer_0[3694] ^ layer_0[254]); 
    assign out[1066] = layer_0[2036]; 
    assign out[1067] = layer_0[525] ^ layer_0[1755]; 
    assign out[1068] = layer_0[2264] & ~layer_0[560]; 
    assign out[1069] = ~(layer_0[3174] & layer_0[3941]); 
    assign out[1070] = layer_0[2052]; 
    assign out[1071] = ~(layer_0[496] ^ layer_0[1707]); 
    assign out[1072] = ~(layer_0[794] ^ layer_0[1382]); 
    assign out[1073] = layer_0[3854]; 
    assign out[1074] = layer_0[2113] & ~layer_0[3066]; 
    assign out[1075] = ~(layer_0[121] | layer_0[2058]); 
    assign out[1076] = layer_0[2818] ^ layer_0[2480]; 
    assign out[1077] = layer_0[29]; 
    assign out[1078] = ~layer_0[1057]; 
    assign out[1079] = ~layer_0[2080]; 
    assign out[1080] = layer_0[2200] & ~layer_0[3159]; 
    assign out[1081] = layer_0[2629] ^ layer_0[1177]; 
    assign out[1082] = ~layer_0[2685]; 
    assign out[1083] = layer_0[3583] ^ layer_0[549]; 
    assign out[1084] = ~(layer_0[1178] ^ layer_0[1964]); 
    assign out[1085] = ~layer_0[2508]; 
    assign out[1086] = layer_0[3315] ^ layer_0[601]; 
    assign out[1087] = ~(layer_0[1624] ^ layer_0[2889]); 
    assign out[1088] = ~(layer_0[2646] | layer_0[2861]); 
    assign out[1089] = layer_0[550]; 
    assign out[1090] = ~(layer_0[3279] ^ layer_0[3114]); 
    assign out[1091] = ~(layer_0[3253] | layer_0[3189]); 
    assign out[1092] = layer_0[1828] ^ layer_0[1110]; 
    assign out[1093] = layer_0[983]; 
    assign out[1094] = ~layer_0[3442]; 
    assign out[1095] = ~layer_0[3427]; 
    assign out[1096] = layer_0[2785]; 
    assign out[1097] = layer_0[2645]; 
    assign out[1098] = ~(layer_0[648] ^ layer_0[3913]); 
    assign out[1099] = ~layer_0[2520]; 
    assign out[1100] = layer_0[1760] & ~layer_0[779]; 
    assign out[1101] = ~layer_0[1208] | (layer_0[1208] & layer_0[3874]); 
    assign out[1102] = layer_0[3706]; 
    assign out[1103] = layer_0[2532]; 
    assign out[1104] = layer_0[2598] & ~layer_0[973]; 
    assign out[1105] = layer_0[3205]; 
    assign out[1106] = ~layer_0[1632]; 
    assign out[1107] = ~(layer_0[3212] | layer_0[2214]); 
    assign out[1108] = ~(layer_0[2503] | layer_0[891]); 
    assign out[1109] = ~layer_0[1955]; 
    assign out[1110] = layer_0[3677] ^ layer_0[1242]; 
    assign out[1111] = ~layer_0[1090]; 
    assign out[1112] = layer_0[268] ^ layer_0[3112]; 
    assign out[1113] = layer_0[259] ^ layer_0[2393]; 
    assign out[1114] = layer_0[2928]; 
    assign out[1115] = layer_0[3868]; 
    assign out[1116] = ~(layer_0[706] ^ layer_0[39]); 
    assign out[1117] = layer_0[17] & ~layer_0[3691]; 
    assign out[1118] = layer_0[375] & layer_0[2038]; 
    assign out[1119] = layer_0[491] & ~layer_0[1432]; 
    assign out[1120] = ~(layer_0[1023] ^ layer_0[1773]); 
    assign out[1121] = layer_0[94] | layer_0[1487]; 
    assign out[1122] = ~layer_0[765]; 
    assign out[1123] = layer_0[675] ^ layer_0[2157]; 
    assign out[1124] = layer_0[2307] ^ layer_0[3451]; 
    assign out[1125] = layer_0[2940]; 
    assign out[1126] = layer_0[3094] & layer_0[430]; 
    assign out[1127] = ~layer_0[1703]; 
    assign out[1128] = layer_0[480]; 
    assign out[1129] = layer_0[882] & ~layer_0[31]; 
    assign out[1130] = ~(layer_0[1256] | layer_0[437]); 
    assign out[1131] = ~(layer_0[1203] ^ layer_0[2403]); 
    assign out[1132] = ~layer_0[1960]; 
    assign out[1133] = ~(layer_0[3025] ^ layer_0[3433]); 
    assign out[1134] = ~layer_0[55]; 
    assign out[1135] = ~(layer_0[3063] ^ layer_0[2912]); 
    assign out[1136] = ~layer_0[2627]; 
    assign out[1137] = ~(layer_0[3339] | layer_0[3716]); 
    assign out[1138] = layer_0[3782] ^ layer_0[2679]; 
    assign out[1139] = ~(layer_0[1002] | layer_0[3921]); 
    assign out[1140] = ~layer_0[1305]; 
    assign out[1141] = ~layer_0[478]; 
    assign out[1142] = layer_0[3898] ^ layer_0[3152]; 
    assign out[1143] = layer_0[2432]; 
    assign out[1144] = ~(layer_0[279] ^ layer_0[2410]); 
    assign out[1145] = layer_0[1746]; 
    assign out[1146] = ~(layer_0[3484] | layer_0[1417]); 
    assign out[1147] = layer_0[2892] & ~layer_0[3690]; 
    assign out[1148] = layer_0[1351] ^ layer_0[1765]; 
    assign out[1149] = ~layer_0[2292]; 
    assign out[1150] = ~(layer_0[1420] ^ layer_0[451]); 
    assign out[1151] = layer_0[2865]; 
    assign out[1152] = ~(layer_0[948] ^ layer_0[1692]); 
    assign out[1153] = layer_0[273] & ~layer_0[209]; 
    assign out[1154] = ~(layer_0[2364] ^ layer_0[755]); 
    assign out[1155] = layer_0[3736] & layer_0[2099]; 
    assign out[1156] = layer_0[502] & ~layer_0[167]; 
    assign out[1157] = layer_0[246] | layer_0[1370]; 
    assign out[1158] = layer_0[754]; 
    assign out[1159] = layer_0[1126] ^ layer_0[2751]; 
    assign out[1160] = layer_0[2585] & ~layer_0[2502]; 
    assign out[1161] = layer_0[3498]; 
    assign out[1162] = ~(layer_0[2358] | layer_0[1211]); 
    assign out[1163] = layer_0[3459] ^ layer_0[3117]; 
    assign out[1164] = ~(layer_0[2711] ^ layer_0[1684]); 
    assign out[1165] = layer_0[3249] ^ layer_0[3366]; 
    assign out[1166] = ~(layer_0[3376] ^ layer_0[3215]); 
    assign out[1167] = layer_0[3170]; 
    assign out[1168] = layer_0[3764] ^ layer_0[139]; 
    assign out[1169] = ~(layer_0[776] & layer_0[3673]); 
    assign out[1170] = ~(layer_0[2570] | layer_0[13]); 
    assign out[1171] = ~layer_0[1955]; 
    assign out[1172] = layer_0[2934] ^ layer_0[101]; 
    assign out[1173] = layer_0[3766] ^ layer_0[1069]; 
    assign out[1174] = ~layer_0[3252]; 
    assign out[1175] = ~(layer_0[3405] ^ layer_0[2578]); 
    assign out[1176] = ~(layer_0[2981] | layer_0[3122]); 
    assign out[1177] = layer_0[22] ^ layer_0[2371]; 
    assign out[1178] = layer_0[2380] & ~layer_0[3958]; 
    assign out[1179] = ~(layer_0[2316] ^ layer_0[3276]); 
    assign out[1180] = layer_0[3083] & ~layer_0[2276]; 
    assign out[1181] = layer_0[1643]; 
    assign out[1182] = layer_0[3222] & layer_0[3573]; 
    assign out[1183] = layer_0[352] & ~layer_0[1987]; 
    assign out[1184] = ~(layer_0[465] ^ layer_0[2389]); 
    assign out[1185] = layer_0[681]; 
    assign out[1186] = ~layer_0[884]; 
    assign out[1187] = ~(layer_0[2902] ^ layer_0[2660]); 
    assign out[1188] = ~layer_0[30]; 
    assign out[1189] = ~(layer_0[2] ^ layer_0[3061]); 
    assign out[1190] = ~(layer_0[3157] ^ layer_0[412]); 
    assign out[1191] = ~(layer_0[452] ^ layer_0[312]); 
    assign out[1192] = ~(layer_0[3870] ^ layer_0[612]); 
    assign out[1193] = layer_0[1036] & layer_0[2717]; 
    assign out[1194] = ~layer_0[2767]; 
    assign out[1195] = layer_0[1940] ^ layer_0[2399]; 
    assign out[1196] = layer_0[1908]; 
    assign out[1197] = ~layer_0[613]; 
    assign out[1198] = ~layer_0[1408]; 
    assign out[1199] = ~(layer_0[2978] | layer_0[3073]); 
    assign out[1200] = layer_0[2915] ^ layer_0[1834]; 
    assign out[1201] = ~layer_0[3211]; 
    assign out[1202] = layer_0[3296] ^ layer_0[2695]; 
    assign out[1203] = ~(layer_0[1798] | layer_0[585]); 
    assign out[1204] = layer_0[957] ^ layer_0[2904]; 
    assign out[1205] = layer_0[770]; 
    assign out[1206] = ~(layer_0[551] & layer_0[248]); 
    assign out[1207] = layer_0[926] & ~layer_0[64]; 
    assign out[1208] = ~layer_0[2971] | (layer_0[1409] & layer_0[2971]); 
    assign out[1209] = layer_0[3003]; 
    assign out[1210] = layer_0[214] ^ layer_0[3732]; 
    assign out[1211] = ~layer_0[447]; 
    assign out[1212] = ~(layer_0[736] ^ layer_0[3737]); 
    assign out[1213] = layer_0[3895]; 
    assign out[1214] = layer_0[1598]; 
    assign out[1215] = layer_0[885] ^ layer_0[2495]; 
    assign out[1216] = layer_0[951]; 
    assign out[1217] = layer_0[3476] & ~layer_0[1438]; 
    assign out[1218] = ~layer_0[2496] | (layer_0[2496] & layer_0[1771]); 
    assign out[1219] = ~layer_0[2672]; 
    assign out[1220] = ~layer_0[115]; 
    assign out[1221] = layer_0[2518] & layer_0[1811]; 
    assign out[1222] = layer_0[57] & ~layer_0[3072]; 
    assign out[1223] = layer_0[1106]; 
    assign out[1224] = layer_0[1319] & layer_0[1453]; 
    assign out[1225] = layer_0[1070] & layer_0[305]; 
    assign out[1226] = ~(layer_0[3204] & layer_0[616]); 
    assign out[1227] = ~(layer_0[217] ^ layer_0[2014]); 
    assign out[1228] = ~layer_0[2637]; 
    assign out[1229] = layer_0[3331]; 
    assign out[1230] = ~layer_0[2460]; 
    assign out[1231] = ~(layer_0[2856] ^ layer_0[737]); 
    assign out[1232] = layer_0[307] ^ layer_0[723]; 
    assign out[1233] = ~layer_0[477]; 
    assign out[1234] = ~(layer_0[3974] ^ layer_0[2297]); 
    assign out[1235] = ~(layer_0[1395] ^ layer_0[2919]); 
    assign out[1236] = layer_0[2185] ^ layer_0[576]; 
    assign out[1237] = ~layer_0[2970]; 
    assign out[1238] = layer_0[3639]; 
    assign out[1239] = ~(layer_0[3491] & layer_0[198]); 
    assign out[1240] = layer_0[62] ^ layer_0[2737]; 
    assign out[1241] = layer_0[2120] ^ layer_0[1060]; 
    assign out[1242] = layer_0[3133] ^ layer_0[939]; 
    assign out[1243] = ~(layer_0[1489] & layer_0[3423]); 
    assign out[1244] = layer_0[1077] ^ layer_0[1045]; 
    assign out[1245] = layer_0[2318] & ~layer_0[1037]; 
    assign out[1246] = layer_0[1606]; 
    assign out[1247] = ~layer_0[3832] | (layer_0[3832] & layer_0[2903]); 
    assign out[1248] = ~layer_0[2485]; 
    assign out[1249] = layer_0[1922] ^ layer_0[3995]; 
    assign out[1250] = ~layer_0[2581]; 
    assign out[1251] = layer_0[25]; 
    assign out[1252] = ~(layer_0[657] | layer_0[247]); 
    assign out[1253] = ~(layer_0[606] | layer_0[927]); 
    assign out[1254] = ~layer_0[1162]; 
    assign out[1255] = layer_0[3715] & ~layer_0[2436]; 
    assign out[1256] = ~(layer_0[2372] ^ layer_0[2510]); 
    assign out[1257] = layer_0[1299] ^ layer_0[669]; 
    assign out[1258] = layer_0[1086] ^ layer_0[2083]; 
    assign out[1259] = ~layer_0[3389]; 
    assign out[1260] = layer_0[1055] | layer_0[2809]; 
    assign out[1261] = ~layer_0[2153]; 
    assign out[1262] = ~layer_0[103] | (layer_0[3785] & layer_0[103]); 
    assign out[1263] = layer_0[2424] & ~layer_0[2924]; 
    assign out[1264] = ~(layer_0[2240] ^ layer_0[528]); 
    assign out[1265] = layer_0[2938]; 
    assign out[1266] = ~(layer_0[2054] & layer_0[3403]); 
    assign out[1267] = ~layer_0[1353]; 
    assign out[1268] = ~layer_0[1329]; 
    assign out[1269] = layer_0[3383] | layer_0[928]; 
    assign out[1270] = ~layer_0[2272]; 
    assign out[1271] = layer_0[1492]; 
    assign out[1272] = ~layer_0[3722] | (layer_0[3957] & layer_0[3722]); 
    assign out[1273] = ~layer_0[3460]; 
    assign out[1274] = ~(layer_0[2523] & layer_0[3208]); 
    assign out[1275] = layer_0[3140]; 
    assign out[1276] = ~layer_0[1147] | (layer_0[1164] & layer_0[1147]); 
    assign out[1277] = layer_0[3892] ^ layer_0[1005]; 
    assign out[1278] = ~layer_0[582]; 
    assign out[1279] = ~layer_0[607]; 
    assign out[1280] = layer_0[3755]; 
    assign out[1281] = layer_0[949] & layer_0[3938]; 
    assign out[1282] = layer_0[600] ^ layer_0[2029]; 
    assign out[1283] = ~(layer_0[2708] ^ layer_0[3455]); 
    assign out[1284] = ~(layer_0[3153] ^ layer_0[3763]); 
    assign out[1285] = ~(layer_0[436] & layer_0[3750]); 
    assign out[1286] = ~layer_0[1582] | (layer_0[1582] & layer_0[2650]); 
    assign out[1287] = ~layer_0[499] | (layer_0[2925] & layer_0[499]); 
    assign out[1288] = layer_0[3685]; 
    assign out[1289] = layer_0[2847] ^ layer_0[1898]; 
    assign out[1290] = ~(layer_0[836] ^ layer_0[2681]); 
    assign out[1291] = ~(layer_0[3246] ^ layer_0[1610]); 
    assign out[1292] = layer_0[3667] ^ layer_0[2395]; 
    assign out[1293] = layer_0[531]; 
    assign out[1294] = layer_0[117] ^ layer_0[653]; 
    assign out[1295] = layer_0[114]; 
    assign out[1296] = layer_0[1630] ^ layer_0[817]; 
    assign out[1297] = layer_0[1501] & layer_0[3501]; 
    assign out[1298] = layer_0[1395]; 
    assign out[1299] = layer_0[1003] & ~layer_0[2051]; 
    assign out[1300] = ~layer_0[3927]; 
    assign out[1301] = ~layer_0[806] | (layer_0[3187] & layer_0[806]); 
    assign out[1302] = ~(layer_0[2884] ^ layer_0[0]); 
    assign out[1303] = layer_0[535] ^ layer_0[1577]; 
    assign out[1304] = layer_0[1346] & ~layer_0[152]; 
    assign out[1305] = ~(layer_0[3128] ^ layer_0[1049]); 
    assign out[1306] = ~(layer_0[810] ^ layer_0[2601]); 
    assign out[1307] = layer_0[3527] ^ layer_0[1206]; 
    assign out[1308] = layer_0[3606]; 
    assign out[1309] = layer_0[1358]; 
    assign out[1310] = layer_0[3421]; 
    assign out[1311] = layer_0[1410]; 
    assign out[1312] = layer_0[2713] ^ layer_0[832]; 
    assign out[1313] = layer_0[628]; 
    assign out[1314] = layer_0[2060]; 
    assign out[1315] = ~(layer_0[1912] ^ layer_0[3040]); 
    assign out[1316] = layer_0[120] & ~layer_0[3535]; 
    assign out[1317] = ~layer_0[1058]; 
    assign out[1318] = layer_0[1482]; 
    assign out[1319] = ~(layer_0[1033] ^ layer_0[1293]); 
    assign out[1320] = ~(layer_0[3797] ^ layer_0[1286]); 
    assign out[1321] = layer_0[3173] ^ layer_0[1454]; 
    assign out[1322] = ~(layer_0[2164] ^ layer_0[3794]); 
    assign out[1323] = ~(layer_0[1118] ^ layer_0[3470]); 
    assign out[1324] = ~layer_0[823] | (layer_0[985] & layer_0[823]); 
    assign out[1325] = layer_0[310] ^ layer_0[3006]; 
    assign out[1326] = ~(layer_0[3646] ^ layer_0[1404]); 
    assign out[1327] = ~layer_0[2107]; 
    assign out[1328] = layer_0[3191]; 
    assign out[1329] = ~layer_0[1669]; 
    assign out[1330] = ~layer_0[3201]; 
    assign out[1331] = ~(layer_0[3334] ^ layer_0[3000]); 
    assign out[1332] = ~layer_0[2152]; 
    assign out[1333] = ~layer_0[3594]; 
    assign out[1334] = layer_0[156]; 
    assign out[1335] = ~(layer_0[2350] ^ layer_0[3815]); 
    assign out[1336] = layer_0[260] & ~layer_0[1693]; 
    assign out[1337] = layer_0[2779]; 
    assign out[1338] = layer_0[2615] & ~layer_0[1238]; 
    assign out[1339] = layer_0[1276]; 
    assign out[1340] = layer_0[2870]; 
    assign out[1341] = layer_0[916]; 
    assign out[1342] = ~(layer_0[2207] ^ layer_0[1136]); 
    assign out[1343] = layer_0[1013]; 
    assign out[1344] = ~layer_0[604] | (layer_0[604] & layer_0[3771]); 
    assign out[1345] = layer_0[2231]; 
    assign out[1346] = layer_0[3370]; 
    assign out[1347] = layer_0[2442]; 
    assign out[1348] = ~(layer_0[266] & layer_0[1028]); 
    assign out[1349] = ~layer_0[1488]; 
    assign out[1350] = ~layer_0[697]; 
    assign out[1351] = ~(layer_0[2920] ^ layer_0[3458]); 
    assign out[1352] = layer_0[1856]; 
    assign out[1353] = layer_0[2735] | layer_0[1318]; 
    assign out[1354] = ~(layer_0[1198] | layer_0[2848]); 
    assign out[1355] = ~(layer_0[1830] ^ layer_0[42]); 
    assign out[1356] = ~(layer_0[3102] & layer_0[2445]); 
    assign out[1357] = layer_0[3733] & ~layer_0[1621]; 
    assign out[1358] = layer_0[3081] ^ layer_0[3486]; 
    assign out[1359] = ~layer_0[2340] | (layer_0[2065] & layer_0[2340]); 
    assign out[1360] = layer_0[3037] & ~layer_0[1507]; 
    assign out[1361] = ~layer_0[2723]; 
    assign out[1362] = layer_0[2554]; 
    assign out[1363] = layer_0[1179]; 
    assign out[1364] = ~(layer_0[1500] ^ layer_0[428]); 
    assign out[1365] = ~layer_0[1853]; 
    assign out[1366] = ~layer_0[1467] | (layer_0[1467] & layer_0[1780]); 
    assign out[1367] = ~(layer_0[1791] & layer_0[1927]); 
    assign out[1368] = layer_0[3565] & ~layer_0[1802]; 
    assign out[1369] = ~(layer_0[2361] ^ layer_0[961]); 
    assign out[1370] = layer_0[664] | layer_0[3027]; 
    assign out[1371] = ~layer_0[1491]; 
    assign out[1372] = layer_0[803] & ~layer_0[3239]; 
    assign out[1373] = layer_0[3397]; 
    assign out[1374] = layer_0[2777]; 
    assign out[1375] = layer_0[3410]; 
    assign out[1376] = ~layer_0[2265] | (layer_0[2977] & layer_0[2265]); 
    assign out[1377] = layer_0[3811]; 
    assign out[1378] = ~layer_0[3062]; 
    assign out[1379] = ~layer_0[2466] | (layer_0[2466] & layer_0[2543]); 
    assign out[1380] = ~layer_0[3444] | (layer_0[3444] & layer_0[1508]); 
    assign out[1381] = layer_0[3580]; 
    assign out[1382] = layer_0[1002]; 
    assign out[1383] = ~(layer_0[448] ^ layer_0[3036]); 
    assign out[1384] = layer_0[1005] ^ layer_0[1942]; 
    assign out[1385] = ~(layer_0[3447] ^ layer_0[1437]); 
    assign out[1386] = layer_0[3339]; 
    assign out[1387] = ~(layer_0[2647] ^ layer_0[536]); 
    assign out[1388] = layer_0[379] & ~layer_0[3247]; 
    assign out[1389] = ~(layer_0[1271] & layer_0[323]); 
    assign out[1390] = layer_0[598] ^ layer_0[1848]; 
    assign out[1391] = layer_0[2703] & layer_0[2150]; 
    assign out[1392] = ~(layer_0[2249] | layer_0[2249]); 
    assign out[1393] = layer_0[2710]; 
    assign out[1394] = ~layer_0[704]; 
    assign out[1395] = layer_0[3364] & ~layer_0[3730]; 
    assign out[1396] = layer_0[238] & layer_0[2692]; 
    assign out[1397] = layer_0[3028] ^ layer_0[792]; 
    assign out[1398] = layer_0[844]; 
    assign out[1399] = layer_0[3355] ^ layer_0[2279]; 
    assign out[1400] = ~(layer_0[590] ^ layer_0[2182]); 
    assign out[1401] = layer_0[3707] | layer_0[137]; 
    assign out[1402] = ~layer_0[2355] | (layer_0[2355] & layer_0[3231]); 
    assign out[1403] = ~(layer_0[1022] ^ layer_0[719]); 
    assign out[1404] = layer_0[3858]; 
    assign out[1405] = layer_0[1982]; 
    assign out[1406] = ~layer_0[2457]; 
    assign out[1407] = ~(layer_0[1687] ^ layer_0[3631]); 
    assign out[1408] = layer_0[2192] ^ layer_0[2505]; 
    assign out[1409] = layer_0[3254]; 
    assign out[1410] = ~layer_0[1074]; 
    assign out[1411] = ~layer_0[660] | (layer_0[49] & layer_0[660]); 
    assign out[1412] = ~layer_0[1557]; 
    assign out[1413] = layer_0[3349] | layer_0[1253]; 
    assign out[1414] = layer_0[1338] ^ layer_0[2370]; 
    assign out[1415] = ~layer_0[2354]; 
    assign out[1416] = layer_0[1336] ^ layer_0[2846]; 
    assign out[1417] = ~layer_0[418]; 
    assign out[1418] = layer_0[596] & layer_0[1174]; 
    assign out[1419] = ~layer_0[645]; 
    assign out[1420] = ~(layer_0[132] ^ layer_0[3700]); 
    assign out[1421] = layer_0[348] ^ layer_0[3305]; 
    assign out[1422] = ~layer_0[864]; 
    assign out[1423] = layer_0[243] & ~layer_0[1255]; 
    assign out[1424] = layer_0[365] & ~layer_0[2241]; 
    assign out[1425] = ~layer_0[492]; 
    assign out[1426] = ~(layer_0[1974] & layer_0[1768]); 
    assign out[1427] = layer_0[1103]; 
    assign out[1428] = ~layer_0[2569]; 
    assign out[1429] = layer_0[2691]; 
    assign out[1430] = layer_0[3997]; 
    assign out[1431] = ~(layer_0[1077] ^ layer_0[1295]); 
    assign out[1432] = layer_0[429]; 
    assign out[1433] = layer_0[75] & ~layer_0[1232]; 
    assign out[1434] = ~layer_0[2089]; 
    assign out[1435] = layer_0[1690] ^ layer_0[725]; 
    assign out[1436] = layer_0[1998]; 
    assign out[1437] = layer_0[762] & layer_0[308]; 
    assign out[1438] = layer_0[3897] ^ layer_0[761]; 
    assign out[1439] = ~(layer_0[168] ^ layer_0[3507]); 
    assign out[1440] = ~(layer_0[1830] ^ layer_0[2729]); 
    assign out[1441] = layer_0[2564]; 
    assign out[1442] = layer_0[3724] ^ layer_0[2843]; 
    assign out[1443] = ~layer_0[3391]; 
    assign out[1444] = ~(layer_0[3144] & layer_0[1689]); 
    assign out[1445] = layer_0[575] & ~layer_0[2188]; 
    assign out[1446] = layer_0[3150]; 
    assign out[1447] = layer_0[3082] & ~layer_0[2754]; 
    assign out[1448] = layer_0[3878] ^ layer_0[177]; 
    assign out[1449] = ~(layer_0[790] ^ layer_0[3281]); 
    assign out[1450] = layer_0[1792] | layer_0[2481]; 
    assign out[1451] = ~(layer_0[3857] & layer_0[619]); 
    assign out[1452] = ~layer_0[3020] | (layer_0[159] & layer_0[3020]); 
    assign out[1453] = ~(layer_0[3575] ^ layer_0[3886]); 
    assign out[1454] = ~(layer_0[1857] ^ layer_0[3668]); 
    assign out[1455] = ~layer_0[56]; 
    assign out[1456] = layer_0[450] & ~layer_0[332]; 
    assign out[1457] = ~(layer_0[2380] | layer_0[3926]); 
    assign out[1458] = layer_0[396]; 
    assign out[1459] = ~(layer_0[1526] ^ layer_0[3684]); 
    assign out[1460] = layer_0[2987] ^ layer_0[2117]; 
    assign out[1461] = layer_0[2084] | layer_0[72]; 
    assign out[1462] = ~(layer_0[3792] ^ layer_0[3934]); 
    assign out[1463] = layer_0[3186] | layer_0[2388]; 
    assign out[1464] = ~(layer_0[2862] ^ layer_0[1561]); 
    assign out[1465] = layer_0[1646] & ~layer_0[2929]; 
    assign out[1466] = layer_0[913]; 
    assign out[1467] = layer_0[1797]; 
    assign out[1468] = ~(layer_0[3980] ^ layer_0[2614]); 
    assign out[1469] = ~layer_0[3515] | (layer_0[3515] & layer_0[986]); 
    assign out[1470] = layer_0[1812]; 
    assign out[1471] = ~layer_0[3505] | (layer_0[1438] & layer_0[3505]); 
    assign out[1472] = ~(layer_0[992] | layer_0[1317]); 
    assign out[1473] = layer_0[1609] ^ layer_0[3975]; 
    assign out[1474] = ~layer_0[1440] | (layer_0[1440] & layer_0[1593]); 
    assign out[1475] = layer_0[2835]; 
    assign out[1476] = ~layer_0[2592]; 
    assign out[1477] = ~layer_0[2147]; 
    assign out[1478] = layer_0[3850] ^ layer_0[370]; 
    assign out[1479] = layer_0[2817] ^ layer_0[759]; 
    assign out[1480] = ~layer_0[3003]; 
    assign out[1481] = layer_0[1631] & ~layer_0[3234]; 
    assign out[1482] = layer_0[567] ^ layer_0[2952]; 
    assign out[1483] = ~(layer_0[3319] ^ layer_0[2568]); 
    assign out[1484] = layer_0[2280] & ~layer_0[670]; 
    assign out[1485] = layer_0[337] ^ layer_0[293]; 
    assign out[1486] = layer_0[3396] ^ layer_0[2434]; 
    assign out[1487] = layer_0[1169] ^ layer_0[2580]; 
    assign out[1488] = layer_0[2501] & ~layer_0[3274]; 
    assign out[1489] = layer_0[3472] ^ layer_0[1633]; 
    assign out[1490] = layer_0[2438] & ~layer_0[183]; 
    assign out[1491] = layer_0[1520] & ~layer_0[3050]; 
    assign out[1492] = ~(layer_0[678] | layer_0[2965]); 
    assign out[1493] = layer_0[1278] ^ layer_0[36]; 
    assign out[1494] = layer_0[3916]; 
    assign out[1495] = ~(layer_0[3225] | layer_0[1936]); 
    assign out[1496] = layer_0[2247] ^ layer_0[1552]; 
    assign out[1497] = layer_0[3008] & ~layer_0[57]; 
    assign out[1498] = layer_0[3626] ^ layer_0[1081]; 
    assign out[1499] = layer_0[1849] ^ layer_0[2329]; 
    assign out[1500] = ~layer_0[1753]; 
    assign out[1501] = ~(layer_0[3553] ^ layer_0[2234]); 
    assign out[1502] = ~layer_0[2000]; 
    assign out[1503] = ~layer_0[2891] | (layer_0[758] & layer_0[2891]); 
    assign out[1504] = layer_0[1085] & ~layer_0[1447]; 
    assign out[1505] = layer_0[377] ^ layer_0[3475]; 
    assign out[1506] = ~(layer_0[2376] & layer_0[2584]); 
    assign out[1507] = layer_0[1997] ^ layer_0[2407]; 
    assign out[1508] = ~(layer_0[3171] ^ layer_0[702]); 
    assign out[1509] = layer_0[3528]; 
    assign out[1510] = layer_0[1085]; 
    assign out[1511] = ~layer_0[3226]; 
    assign out[1512] = layer_0[81] & layer_0[219]; 
    assign out[1513] = ~layer_0[1876]; 
    assign out[1514] = ~(layer_0[1048] ^ layer_0[2797]); 
    assign out[1515] = ~(layer_0[3807] ^ layer_0[2377]); 
    assign out[1516] = layer_0[1001]; 
    assign out[1517] = ~layer_0[3462]; 
    assign out[1518] = ~layer_0[1400]; 
    assign out[1519] = ~layer_0[124]; 
    assign out[1520] = ~layer_0[733] | (layer_0[1021] & layer_0[733]); 
    assign out[1521] = ~(layer_0[1046] ^ layer_0[3340]); 
    assign out[1522] = layer_0[3196] ^ layer_0[1130]; 
    assign out[1523] = layer_0[1331]; 
    assign out[1524] = ~(layer_0[3394] ^ layer_0[1080]); 
    assign out[1525] = layer_0[2165] ^ layer_0[838]; 
    assign out[1526] = layer_0[1487] & layer_0[1894]; 
    assign out[1527] = layer_0[2816] ^ layer_0[2441]; 
    assign out[1528] = ~(layer_0[1771] | layer_0[1225]); 
    assign out[1529] = ~layer_0[3304] | (layer_0[3714] & layer_0[3304]); 
    assign out[1530] = ~(layer_0[345] ^ layer_0[3308]); 
    assign out[1531] = layer_0[2374] & ~layer_0[3978]; 
    assign out[1532] = layer_0[1641] & ~layer_0[1321]; 
    assign out[1533] = layer_0[472] ^ layer_0[1973]; 
    assign out[1534] = layer_0[724]; 
    assign out[1535] = layer_0[505]; 
    assign out[1536] = ~layer_0[2367]; 
    assign out[1537] = ~layer_0[288]; 
    assign out[1538] = layer_0[815] ^ layer_0[3791]; 
    assign out[1539] = ~layer_0[2319]; 
    assign out[1540] = layer_0[845] ^ layer_0[3069]; 
    assign out[1541] = ~layer_0[630]; 
    assign out[1542] = layer_0[1326] ^ layer_0[2255]; 
    assign out[1543] = layer_0[525]; 
    assign out[1544] = layer_0[714] & layer_0[1383]; 
    assign out[1545] = layer_0[3026] ^ layer_0[3560]; 
    assign out[1546] = layer_0[2743] & ~layer_0[2997]; 
    assign out[1547] = layer_0[3306] ^ layer_0[2741]; 
    assign out[1548] = ~(layer_0[3273] | layer_0[1924]); 
    assign out[1549] = ~layer_0[3798]; 
    assign out[1550] = layer_0[1503] & ~layer_0[893]; 
    assign out[1551] = ~layer_0[397]; 
    assign out[1552] = layer_0[1890]; 
    assign out[1553] = ~(layer_0[2531] | layer_0[2296]); 
    assign out[1554] = ~(layer_0[2854] & layer_0[232]); 
    assign out[1555] = layer_0[3601] & ~layer_0[2828]; 
    assign out[1556] = layer_0[757] & ~layer_0[3413]; 
    assign out[1557] = ~layer_0[514]; 
    assign out[1558] = layer_0[3231]; 
    assign out[1559] = ~(layer_0[2020] ^ layer_0[3863]); 
    assign out[1560] = ~layer_0[3210]; 
    assign out[1561] = ~(layer_0[1295] ^ layer_0[483]); 
    assign out[1562] = ~layer_0[633]; 
    assign out[1563] = layer_0[3780] & layer_0[90]; 
    assign out[1564] = layer_0[1028] & layer_0[271]; 
    assign out[1565] = ~(layer_0[3504] | layer_0[2115]); 
    assign out[1566] = layer_0[3682]; 
    assign out[1567] = layer_0[705] ^ layer_0[223]; 
    assign out[1568] = layer_0[3298]; 
    assign out[1569] = layer_0[1303]; 
    assign out[1570] = layer_0[501] ^ layer_0[2181]; 
    assign out[1571] = layer_0[1992] ^ layer_0[3322]; 
    assign out[1572] = ~(layer_0[3820] ^ layer_0[448]); 
    assign out[1573] = ~layer_0[2516]; 
    assign out[1574] = layer_0[3513]; 
    assign out[1575] = ~layer_0[3742]; 
    assign out[1576] = layer_0[2879]; 
    assign out[1577] = layer_0[2528]; 
    assign out[1578] = ~(layer_0[937] ^ layer_0[3437]); 
    assign out[1579] = layer_0[2308] ^ layer_0[3384]; 
    assign out[1580] = ~(layer_0[2608] | layer_0[1223]); 
    assign out[1581] = ~layer_0[837] | (layer_0[3960] & layer_0[837]); 
    assign out[1582] = layer_0[3282] & ~layer_0[3559]; 
    assign out[1583] = ~layer_0[1581]; 
    assign out[1584] = layer_0[652]; 
    assign out[1585] = layer_0[2403]; 
    assign out[1586] = layer_0[1009] & layer_0[2382]; 
    assign out[1587] = layer_0[2664] ^ layer_0[2213]; 
    assign out[1588] = ~(layer_0[1608] ^ layer_0[3045]); 
    assign out[1589] = layer_0[3463] | layer_0[1051]; 
    assign out[1590] = layer_0[178]; 
    assign out[1591] = layer_0[1146] & layer_0[3300]; 
    assign out[1592] = layer_0[2304] | layer_0[612]; 
    assign out[1593] = layer_0[1541] & ~layer_0[640]; 
    assign out[1594] = ~(layer_0[545] ^ layer_0[1356]); 
    assign out[1595] = ~layer_0[1416]; 
    assign out[1596] = ~(layer_0[3628] | layer_0[2560]); 
    assign out[1597] = ~layer_0[1043] | (layer_0[1043] & layer_0[3581]); 
    assign out[1598] = ~(layer_0[1648] ^ layer_0[3786]); 
    assign out[1599] = layer_0[1584] & layer_0[2842]; 
    assign out[1600] = layer_0[2756] & ~layer_0[1845]; 
    assign out[1601] = layer_0[46] ^ layer_0[3866]; 
    assign out[1602] = ~(layer_0[1270] ^ layer_0[2339]); 
    assign out[1603] = layer_0[2452] & layer_0[3043]; 
    assign out[1604] = ~layer_0[3903]; 
    assign out[1605] = ~layer_0[3697]; 
    assign out[1606] = ~(layer_0[3108] ^ layer_0[3610]); 
    assign out[1607] = layer_0[2095]; 
    assign out[1608] = layer_0[2024]; 
    assign out[1609] = layer_0[1545] & ~layer_0[2379]; 
    assign out[1610] = layer_0[764] & ~layer_0[2167]; 
    assign out[1611] = ~layer_0[3520]; 
    assign out[1612] = ~layer_0[3068] | (layer_0[1245] & layer_0[3068]); 
    assign out[1613] = ~layer_0[2469]; 
    assign out[1614] = ~layer_0[146]; 
    assign out[1615] = ~layer_0[873]; 
    assign out[1616] = layer_0[1525] & layer_0[70]; 
    assign out[1617] = layer_0[634]; 
    assign out[1618] = ~(layer_0[398] ^ layer_0[1493]); 
    assign out[1619] = ~(layer_0[2475] ^ layer_0[299]); 
    assign out[1620] = layer_0[590] & ~layer_0[2911]; 
    assign out[1621] = ~(layer_0[3287] ^ layer_0[2449]); 
    assign out[1622] = layer_0[741] ^ layer_0[3248]; 
    assign out[1623] = ~layer_0[835]; 
    assign out[1624] = layer_0[2597]; 
    assign out[1625] = ~(layer_0[1525] ^ layer_0[1257]); 
    assign out[1626] = ~(layer_0[3980] ^ layer_0[2424]); 
    assign out[1627] = ~layer_0[2628]; 
    assign out[1628] = layer_0[3190] ^ layer_0[321]; 
    assign out[1629] = ~(layer_0[2813] ^ layer_0[171]); 
    assign out[1630] = layer_0[824] & layer_0[3385]; 
    assign out[1631] = layer_0[3536] & layer_0[666]; 
    assign out[1632] = ~layer_0[626]; 
    assign out[1633] = layer_0[3358] ^ layer_0[1391]; 
    assign out[1634] = ~(layer_0[644] | layer_0[3279]); 
    assign out[1635] = layer_0[2156] & ~layer_0[1321]; 
    assign out[1636] = ~layer_0[1953]; 
    assign out[1637] = ~layer_0[3312]; 
    assign out[1638] = layer_0[2585] & ~layer_0[1556]; 
    assign out[1639] = layer_0[346] ^ layer_0[2352]; 
    assign out[1640] = ~(layer_0[3012] ^ layer_0[1111]); 
    assign out[1641] = layer_0[2137] & ~layer_0[414]; 
    assign out[1642] = ~layer_0[529]; 
    assign out[1643] = layer_0[1497] & layer_0[2071]; 
    assign out[1644] = layer_0[2934] & ~layer_0[2726]; 
    assign out[1645] = ~(layer_0[3172] | layer_0[2351]); 
    assign out[1646] = layer_0[807]; 
    assign out[1647] = layer_0[2950] ^ layer_0[682]; 
    assign out[1648] = ~layer_0[1788] | (layer_0[1919] & layer_0[1788]); 
    assign out[1649] = layer_0[1382] & ~layer_0[736]; 
    assign out[1650] = ~(layer_0[47] | layer_0[1496]); 
    assign out[1651] = ~(layer_0[3187] & layer_0[404]); 
    assign out[1652] = ~layer_0[2489]; 
    assign out[1653] = layer_0[874] ^ layer_0[615]; 
    assign out[1654] = layer_0[1139] & layer_0[2027]; 
    assign out[1655] = ~(layer_0[1939] ^ layer_0[886]); 
    assign out[1656] = layer_0[2610] & ~layer_0[2050]; 
    assign out[1657] = ~layer_0[3683] | (layer_0[3683] & layer_0[3617]); 
    assign out[1658] = ~(layer_0[470] | layer_0[296]); 
    assign out[1659] = layer_0[334] & ~layer_0[955]; 
    assign out[1660] = layer_0[3572] & layer_0[1936]; 
    assign out[1661] = ~(layer_0[2956] ^ layer_0[3328]); 
    assign out[1662] = ~layer_0[1859] | (layer_0[1872] & layer_0[1859]); 
    assign out[1663] = ~layer_0[3531]; 
    assign out[1664] = ~layer_0[1766] | (layer_0[309] & layer_0[1766]); 
    assign out[1665] = ~(layer_0[357] | layer_0[2419]); 
    assign out[1666] = layer_0[1879]; 
    assign out[1667] = ~layer_0[2154]; 
    assign out[1668] = layer_0[1031]; 
    assign out[1669] = layer_0[1712] & ~layer_0[1754]; 
    assign out[1670] = ~(layer_0[2313] | layer_0[1112]); 
    assign out[1671] = ~(layer_0[1579] | layer_0[2701]); 
    assign out[1672] = layer_0[2321] ^ layer_0[2008]; 
    assign out[1673] = ~layer_0[1576]; 
    assign out[1674] = layer_0[1719]; 
    assign out[1675] = ~(layer_0[3086] ^ layer_0[2776]); 
    assign out[1676] = layer_0[3555] & ~layer_0[2138]; 
    assign out[1677] = layer_0[785] & ~layer_0[3199]; 
    assign out[1678] = ~(layer_0[2013] ^ layer_0[3005]); 
    assign out[1679] = ~(layer_0[866] | layer_0[2763]); 
    assign out[1680] = layer_0[1068] ^ layer_0[3278]; 
    assign out[1681] = ~(layer_0[3213] ^ layer_0[2954]); 
    assign out[1682] = ~(layer_0[2805] ^ layer_0[2194]); 
    assign out[1683] = ~(layer_0[982] | layer_0[786]); 
    assign out[1684] = ~layer_0[1304]; 
    assign out[1685] = ~(layer_0[3981] ^ layer_0[319]); 
    assign out[1686] = layer_0[3395]; 
    assign out[1687] = layer_0[959] ^ layer_0[21]; 
    assign out[1688] = ~(layer_0[3642] ^ layer_0[860]); 
    assign out[1689] = ~(layer_0[1272] ^ layer_0[63]); 
    assign out[1690] = ~layer_0[359]; 
    assign out[1691] = ~(layer_0[1450] ^ layer_0[1347]); 
    assign out[1692] = layer_0[3453] & ~layer_0[1341]; 
    assign out[1693] = ~layer_0[2881]; 
    assign out[1694] = ~layer_0[1875]; 
    assign out[1695] = ~(layer_0[328] ^ layer_0[3836]); 
    assign out[1696] = ~layer_0[335]; 
    assign out[1697] = layer_0[2988] & ~layer_0[1035]; 
    assign out[1698] = layer_0[380] ^ layer_0[182]; 
    assign out[1699] = ~layer_0[1308]; 
    assign out[1700] = layer_0[457] & ~layer_0[1089]; 
    assign out[1701] = layer_0[413] & ~layer_0[3161]; 
    assign out[1702] = layer_0[3206] ^ layer_0[1808]; 
    assign out[1703] = ~(layer_0[1724] | layer_0[597]); 
    assign out[1704] = layer_0[3537] ^ layer_0[2472]; 
    assign out[1705] = ~(layer_0[1000] & layer_0[3826]); 
    assign out[1706] = ~layer_0[830]; 
    assign out[1707] = ~(layer_0[344] & layer_0[3589]); 
    assign out[1708] = ~(layer_0[1296] ^ layer_0[516]); 
    assign out[1709] = layer_0[2811]; 
    assign out[1710] = layer_0[629] & layer_0[1054]; 
    assign out[1711] = ~(layer_0[1389] ^ layer_0[2010]); 
    assign out[1712] = layer_0[3435] & ~layer_0[2779]; 
    assign out[1713] = ~(layer_0[1234] ^ layer_0[92]); 
    assign out[1714] = layer_0[2474] ^ layer_0[1934]; 
    assign out[1715] = ~layer_0[3686]; 
    assign out[1716] = ~layer_0[2028] | (layer_0[2028] & layer_0[1730]); 
    assign out[1717] = layer_0[2844] & ~layer_0[3911]; 
    assign out[1718] = ~layer_0[3404]; 
    assign out[1719] = ~layer_0[914]; 
    assign out[1720] = ~layer_0[2726] | (layer_0[2478] & layer_0[2726]); 
    assign out[1721] = layer_0[3831]; 
    assign out[1722] = ~layer_0[804] | (layer_0[804] & layer_0[3213]); 
    assign out[1723] = ~layer_0[2914]; 
    assign out[1724] = ~(layer_0[3158] | layer_0[2868]); 
    assign out[1725] = ~layer_0[3378]; 
    assign out[1726] = layer_0[2838] & ~layer_0[3527]; 
    assign out[1727] = layer_0[1405] ^ layer_0[2171]; 
    assign out[1728] = ~layer_0[3543]; 
    assign out[1729] = layer_0[3390] ^ layer_0[3752]; 
    assign out[1730] = layer_0[2030] & ~layer_0[3494]; 
    assign out[1731] = layer_0[513] & ~layer_0[3021]; 
    assign out[1732] = layer_0[1883]; 
    assign out[1733] = ~layer_0[1469]; 
    assign out[1734] = layer_0[121] ^ layer_0[1505]; 
    assign out[1735] = ~(layer_0[1569] ^ layer_0[2130]); 
    assign out[1736] = layer_0[909] ^ layer_0[143]; 
    assign out[1737] = ~layer_0[949]; 
    assign out[1738] = ~(layer_0[3889] ^ layer_0[2956]); 
    assign out[1739] = layer_0[1971] ^ layer_0[1195]; 
    assign out[1740] = ~(layer_0[2479] | layer_0[783]); 
    assign out[1741] = ~layer_0[2857] | (layer_0[2857] & layer_0[3227]); 
    assign out[1742] = layer_0[2640]; 
    assign out[1743] = ~layer_0[1306]; 
    assign out[1744] = layer_0[878] & ~layer_0[240]; 
    assign out[1745] = ~(layer_0[3934] ^ layer_0[3796]); 
    assign out[1746] = layer_0[2202] ^ layer_0[556]; 
    assign out[1747] = ~(layer_0[3078] & layer_0[1466]); 
    assign out[1748] = layer_0[3419] ^ layer_0[2332]; 
    assign out[1749] = ~(layer_0[730] ^ layer_0[2253]); 
    assign out[1750] = ~(layer_0[176] ^ layer_0[1523]); 
    assign out[1751] = layer_0[145] & ~layer_0[2325]; 
    assign out[1752] = layer_0[530] & ~layer_0[917]; 
    assign out[1753] = ~(layer_0[3620] | layer_0[2571]); 
    assign out[1754] = ~layer_0[1319]; 
    assign out[1755] = ~(layer_0[2512] & layer_0[3817]); 
    assign out[1756] = ~layer_0[3029] | (layer_0[1623] & layer_0[3029]); 
    assign out[1757] = layer_0[1327] & ~layer_0[972]; 
    assign out[1758] = ~(layer_0[1749] ^ layer_0[97]); 
    assign out[1759] = ~(layer_0[3687] ^ layer_0[504]); 
    assign out[1760] = layer_0[227] ^ layer_0[2183]; 
    assign out[1761] = layer_0[1345] ^ layer_0[1555]; 
    assign out[1762] = layer_0[1043] ^ layer_0[1877]; 
    assign out[1763] = ~(layer_0[1279] ^ layer_0[663]); 
    assign out[1764] = layer_0[631] ^ layer_0[3700]; 
    assign out[1765] = ~layer_0[3999]; 
    assign out[1766] = layer_0[3939]; 
    assign out[1767] = layer_0[820] & ~layer_0[3711]; 
    assign out[1768] = ~layer_0[1160]; 
    assign out[1769] = ~(layer_0[3264] ^ layer_0[1839]); 
    assign out[1770] = layer_0[1369] ^ layer_0[1502]; 
    assign out[1771] = ~(layer_0[1323] ^ layer_0[42]); 
    assign out[1772] = ~(layer_0[2778] | layer_0[2328]); 
    assign out[1773] = layer_0[3762]; 
    assign out[1774] = ~layer_0[2995] | (layer_0[2867] & layer_0[2995]); 
    assign out[1775] = layer_0[1644]; 
    assign out[1776] = layer_0[1399] ^ layer_0[2909]; 
    assign out[1777] = ~(layer_0[1138] | layer_0[2560]); 
    assign out[1778] = layer_0[2832]; 
    assign out[1779] = layer_0[1828] & layer_0[2871]; 
    assign out[1780] = layer_0[2926] ^ layer_0[771]; 
    assign out[1781] = ~(layer_0[2583] ^ layer_0[1667]); 
    assign out[1782] = ~(layer_0[2351] ^ layer_0[414]); 
    assign out[1783] = layer_0[456] & ~layer_0[3575]; 
    assign out[1784] = layer_0[843] ^ layer_0[143]; 
    assign out[1785] = layer_0[2263] ^ layer_0[613]; 
    assign out[1786] = layer_0[1650] & layer_0[3949]; 
    assign out[1787] = layer_0[1430] & ~layer_0[746]; 
    assign out[1788] = layer_0[2328]; 
    assign out[1789] = layer_0[3725] & layer_0[467]; 
    assign out[1790] = layer_0[3918] ^ layer_0[1190]; 
    assign out[1791] = ~(layer_0[3163] ^ layer_0[1628]); 
    assign out[1792] = ~(layer_0[3692] ^ layer_0[294]); 
    assign out[1793] = ~(layer_0[808] | layer_0[3766]); 
    assign out[1794] = ~layer_0[2243]; 
    assign out[1795] = layer_0[1350] | layer_0[113]; 
    assign out[1796] = ~(layer_0[1905] ^ layer_0[3947]); 
    assign out[1797] = ~(layer_0[1461] ^ layer_0[3290]); 
    assign out[1798] = ~(layer_0[495] | layer_0[251]); 
    assign out[1799] = layer_0[1354]; 
    assign out[1800] = layer_0[1282] & ~layer_0[772]; 
    assign out[1801] = ~(layer_0[2394] | layer_0[1518]); 
    assign out[1802] = ~(layer_0[1580] ^ layer_0[2731]); 
    assign out[1803] = ~layer_0[2527]; 
    assign out[1804] = layer_0[1277]; 
    assign out[1805] = layer_0[2707] & ~layer_0[958]; 
    assign out[1806] = layer_0[2952] & ~layer_0[61]; 
    assign out[1807] = layer_0[2162] & ~layer_0[2543]; 
    assign out[1808] = layer_0[2218]; 
    assign out[1809] = ~layer_0[2572] | (layer_0[2572] & layer_0[3728]); 
    assign out[1810] = ~(layer_0[1785] ^ layer_0[2384]); 
    assign out[1811] = layer_0[3262] ^ layer_0[3490]; 
    assign out[1812] = ~layer_0[20]; 
    assign out[1813] = ~(layer_0[1063] ^ layer_0[3452]); 
    assign out[1814] = layer_0[2287] & ~layer_0[719]; 
    assign out[1815] = ~layer_0[411]; 
    assign out[1816] = ~(layer_0[1266] ^ layer_0[441]); 
    assign out[1817] = ~layer_0[3956]; 
    assign out[1818] = layer_0[3987] ^ layer_0[2426]; 
    assign out[1819] = layer_0[1030]; 
    assign out[1820] = ~layer_0[1824]; 
    assign out[1821] = ~(layer_0[2033] | layer_0[2391]); 
    assign out[1822] = layer_0[1108] ^ layer_0[3717]; 
    assign out[1823] = ~layer_0[3937] | (layer_0[971] & layer_0[3937]); 
    assign out[1824] = layer_0[2239] & layer_0[3124]; 
    assign out[1825] = layer_0[1869]; 
    assign out[1826] = layer_0[2778] ^ layer_0[2624]; 
    assign out[1827] = layer_0[2118] ^ layer_0[457]; 
    assign out[1828] = layer_0[449]; 
    assign out[1829] = ~(layer_0[2989] | layer_0[3874]); 
    assign out[1830] = layer_0[2158] & layer_0[3706]; 
    assign out[1831] = ~layer_0[14]; 
    assign out[1832] = ~(layer_0[2286] ^ layer_0[2784]); 
    assign out[1833] = layer_0[2254] & layer_0[2353]; 
    assign out[1834] = ~(layer_0[18] & layer_0[3076]); 
    assign out[1835] = layer_0[751] & ~layer_0[1038]; 
    assign out[1836] = ~(layer_0[3799] | layer_0[1142]); 
    assign out[1837] = layer_0[2248]; 
    assign out[1838] = layer_0[877] & ~layer_0[1673]; 
    assign out[1839] = layer_0[3523]; 
    assign out[1840] = layer_0[3856] & ~layer_0[2476]; 
    assign out[1841] = layer_0[2257]; 
    assign out[1842] = ~(layer_0[3452] ^ layer_0[880]); 
    assign out[1843] = ~layer_0[1743] | (layer_0[1743] & layer_0[1311]); 
    assign out[1844] = ~(layer_0[614] ^ layer_0[2936]); 
    assign out[1845] = layer_0[3653] & ~layer_0[2657]; 
    assign out[1846] = ~(layer_0[1659] ^ layer_0[173]); 
    assign out[1847] = ~layer_0[6] | (layer_0[6] & layer_0[3809]); 
    assign out[1848] = ~(layer_0[3756] ^ layer_0[977]); 
    assign out[1849] = layer_0[3221] | layer_0[3910]; 
    assign out[1850] = layer_0[2245]; 
    assign out[1851] = ~(layer_0[914] ^ layer_0[2224]); 
    assign out[1852] = ~(layer_0[3293] ^ layer_0[1626]); 
    assign out[1853] = ~layer_0[2123] | (layer_0[2869] & layer_0[2123]); 
    assign out[1854] = layer_0[940] | layer_0[1966]; 
    assign out[1855] = layer_0[1559] & layer_0[3949]; 
    assign out[1856] = layer_0[2044] & ~layer_0[3027]; 
    assign out[1857] = layer_0[3194] & ~layer_0[1224]; 
    assign out[1858] = ~layer_0[507]; 
    assign out[1859] = layer_0[1869]; 
    assign out[1860] = ~(layer_0[2841] ^ layer_0[2320]); 
    assign out[1861] = layer_0[1426] & ~layer_0[2298]; 
    assign out[1862] = layer_0[3582] & ~layer_0[754]; 
    assign out[1863] = layer_0[599] & ~layer_0[2208]; 
    assign out[1864] = layer_0[3574] ^ layer_0[434]; 
    assign out[1865] = layer_0[3313] & ~layer_0[61]; 
    assign out[1866] = layer_0[163] & layer_0[1941]; 
    assign out[1867] = layer_0[3739] & ~layer_0[598]; 
    assign out[1868] = layer_0[978] & ~layer_0[1549]; 
    assign out[1869] = ~layer_0[2943] | (layer_0[2943] & layer_0[2819]); 
    assign out[1870] = ~(layer_0[3286] ^ layer_0[2648]); 
    assign out[1871] = layer_0[883] ^ layer_0[1113]; 
    assign out[1872] = layer_0[674] & ~layer_0[1083]; 
    assign out[1873] = ~(layer_0[989] ^ layer_0[2719]); 
    assign out[1874] = layer_0[2807] & layer_0[1468]; 
    assign out[1875] = layer_0[146] & ~layer_0[3042]; 
    assign out[1876] = ~(layer_0[2591] ^ layer_0[2755]); 
    assign out[1877] = layer_0[1027]; 
    assign out[1878] = layer_0[780]; 
    assign out[1879] = layer_0[65] ^ layer_0[2135]; 
    assign out[1880] = ~(layer_0[341] ^ layer_0[3465]); 
    assign out[1881] = layer_0[3804] & ~layer_0[3802]; 
    assign out[1882] = ~(layer_0[3428] ^ layer_0[3162]); 
    assign out[1883] = layer_0[2439]; 
    assign out[1884] = ~(layer_0[1767] | layer_0[2064]); 
    assign out[1885] = ~(layer_0[3541] ^ layer_0[35]); 
    assign out[1886] = ~(layer_0[3740] | layer_0[1268]); 
    assign out[1887] = ~(layer_0[2626] ^ layer_0[3569]); 
    assign out[1888] = ~(layer_0[2860] | layer_0[2907]); 
    assign out[1889] = ~layer_0[1978]; 
    assign out[1890] = layer_0[3857] & ~layer_0[2081]; 
    assign out[1891] = ~(layer_0[2122] | layer_0[2976]); 
    assign out[1892] = ~(layer_0[882] | layer_0[3660]); 
    assign out[1893] = layer_0[3867] ^ layer_0[2177]; 
    assign out[1894] = layer_0[3347] ^ layer_0[3558]; 
    assign out[1895] = ~layer_0[3626]; 
    assign out[1896] = layer_0[2463] & layer_0[1481]; 
    assign out[1897] = layer_0[162] | layer_0[233]; 
    assign out[1898] = ~(layer_0[141] ^ layer_0[2392]); 
    assign out[1899] = layer_0[813] ^ layer_0[3571]; 
    assign out[1900] = ~(layer_0[710] ^ layer_0[2786]); 
    assign out[1901] = layer_0[3344] ^ layer_0[876]; 
    assign out[1902] = layer_0[3482] ^ layer_0[580]; 
    assign out[1903] = ~(layer_0[3160] ^ layer_0[3698]); 
    assign out[1904] = ~layer_0[2942]; 
    assign out[1905] = ~(layer_0[1990] ^ layer_0[2233]); 
    assign out[1906] = layer_0[3188] ^ layer_0[1315]; 
    assign out[1907] = ~(layer_0[1697] ^ layer_0[141]); 
    assign out[1908] = ~(layer_0[988] ^ layer_0[1733]); 
    assign out[1909] = layer_0[1153]; 
    assign out[1910] = layer_0[879] ^ layer_0[41]; 
    assign out[1911] = ~layer_0[2206]; 
    assign out[1912] = ~(layer_0[3977] | layer_0[2062]); 
    assign out[1913] = layer_0[468] & ~layer_0[2360]; 
    assign out[1914] = layer_0[395] ^ layer_0[1256]; 
    assign out[1915] = layer_0[2938]; 
    assign out[1916] = layer_0[1131] ^ layer_0[2720]; 
    assign out[1917] = layer_0[3506] ^ layer_0[2346]; 
    assign out[1918] = ~(layer_0[3765] ^ layer_0[2874]); 
    assign out[1919] = ~(layer_0[3846] ^ layer_0[1625]); 
    assign out[1920] = ~(layer_0[2170] ^ layer_0[3608]); 
    assign out[1921] = ~(layer_0[515] ^ layer_0[1971]); 
    assign out[1922] = layer_0[1404] & ~layer_0[1837]; 
    assign out[1923] = layer_0[2176] ^ layer_0[3539]; 
    assign out[1924] = ~layer_0[829]; 
    assign out[1925] = layer_0[1537] & ~layer_0[218]; 
    assign out[1926] = ~(layer_0[10] ^ layer_0[1320]); 
    assign out[1927] = layer_0[2139]; 
    assign out[1928] = layer_0[3609]; 
    assign out[1929] = ~(layer_0[3417] ^ layer_0[594]); 
    assign out[1930] = ~(layer_0[1886] ^ layer_0[1107]); 
    assign out[1931] = ~(layer_0[853] | layer_0[1340]); 
    assign out[1932] = ~layer_0[3218]; 
    assign out[1933] = layer_0[1784] ^ layer_0[3765]; 
    assign out[1934] = ~(layer_0[742] ^ layer_0[1834]); 
    assign out[1935] = ~(layer_0[119] | layer_0[991]); 
    assign out[1936] = ~layer_0[3059]; 
    assign out[1937] = ~(layer_0[798] ^ layer_0[743]); 
    assign out[1938] = ~(layer_0[1356] ^ layer_0[995]); 
    assign out[1939] = ~(layer_0[1524] | layer_0[2484]); 
    assign out[1940] = ~layer_0[1472] | (layer_0[1472] & layer_0[3753]); 
    assign out[1941] = layer_0[3777] & ~layer_0[2555]; 
    assign out[1942] = ~layer_0[3644] | (layer_0[3644] & layer_0[3611]); 
    assign out[1943] = layer_0[3054] & layer_0[2582]; 
    assign out[1944] = layer_0[2138]; 
    assign out[1945] = ~layer_0[1748]; 
    assign out[1946] = layer_0[2546] ^ layer_0[1294]; 
    assign out[1947] = layer_0[3712] ^ layer_0[2563]; 
    assign out[1948] = ~layer_0[1543]; 
    assign out[1949] = layer_0[2774]; 
    assign out[1950] = layer_0[3948] ^ layer_0[1388]; 
    assign out[1951] = layer_0[1242]; 
    assign out[1952] = ~(layer_0[775] ^ layer_0[771]); 
    assign out[1953] = ~(layer_0[1484] ^ layer_0[3154]); 
    assign out[1954] = ~layer_0[1899] | (layer_0[1899] & layer_0[1162]); 
    assign out[1955] = layer_0[3709] & layer_0[3609]; 
    assign out[1956] = layer_0[3209]; 
    assign out[1957] = layer_0[1260]; 
    assign out[1958] = layer_0[151] ^ layer_0[1948]; 
    assign out[1959] = ~(layer_0[3919] ^ layer_0[2025]); 
    assign out[1960] = ~(layer_0[1723] ^ layer_0[1903]); 
    assign out[1961] = layer_0[1670] & ~layer_0[3236]; 
    assign out[1962] = layer_0[3641] & ~layer_0[3023]; 
    assign out[1963] = ~layer_0[1415]; 
    assign out[1964] = layer_0[2671] ^ layer_0[3621]; 
    assign out[1965] = layer_0[1597] ^ layer_0[2836]; 
    assign out[1966] = ~layer_0[3499]; 
    assign out[1967] = layer_0[1533]; 
    assign out[1968] = layer_0[1448] & ~layer_0[3970]; 
    assign out[1969] = ~layer_0[1812]; 
    assign out[1970] = ~(layer_0[2653] ^ layer_0[3496]); 
    assign out[1971] = ~layer_0[778]; 
    assign out[1972] = ~(layer_0[1882] | layer_0[1301]); 
    assign out[1973] = ~(layer_0[658] ^ layer_0[1744]); 
    assign out[1974] = layer_0[673] ^ layer_0[1386]; 
    assign out[1975] = ~(layer_0[3179] ^ layer_0[301]); 
    assign out[1976] = layer_0[1505] ^ layer_0[1127]; 
    assign out[1977] = layer_0[3607] & ~layer_0[1587]; 
    assign out[1978] = layer_0[687] ^ layer_0[1207]; 
    assign out[1979] = layer_0[2344]; 
    assign out[1980] = ~layer_0[541]; 
    assign out[1981] = layer_0[2369] ^ layer_0[3013]; 
    assign out[1982] = layer_0[3373]; 
    assign out[1983] = layer_0[3] & ~layer_0[872]; 
    assign out[1984] = ~(layer_0[2787] ^ layer_0[3873]); 
    assign out[1985] = ~(layer_0[3469] ^ layer_0[2837]); 
    assign out[1986] = layer_0[2428] ^ layer_0[2097]; 
    assign out[1987] = ~(layer_0[3207] ^ layer_0[37]); 
    assign out[1988] = layer_0[2462]; 
    assign out[1989] = ~(layer_0[3776] ^ layer_0[2872]); 
    assign out[1990] = layer_0[1627] ^ layer_0[1023]; 
    assign out[1991] = ~layer_0[2219]; 
    assign out[1992] = ~(layer_0[2941] ^ layer_0[180]); 
    assign out[1993] = ~layer_0[469]; 
    assign out[1994] = layer_0[2950]; 
    assign out[1995] = layer_0[3779] & ~layer_0[1729]; 
    assign out[1996] = layer_0[336] & layer_0[3654]; 
    assign out[1997] = layer_0[2810] | layer_0[3584]; 
    assign out[1998] = ~layer_0[997]; 
    assign out[1999] = ~(layer_0[2677] ^ layer_0[2878]); 
    assign out[2000] = layer_0[2586] | layer_0[1466]; 
    assign out[2001] = layer_0[3111] & layer_0[1246]; 
    assign out[2002] = ~(layer_0[900] ^ layer_0[1290]); 
    assign out[2003] = ~(layer_0[172] ^ layer_0[2266]); 
    assign out[2004] = ~layer_0[2698] | (layer_0[2698] & layer_0[2819]); 
    assign out[2005] = ~(layer_0[1612] ^ layer_0[387]); 
    assign out[2006] = ~(layer_0[1705] ^ layer_0[2705]); 
    assign out[2007] = layer_0[2335] ^ layer_0[2134]; 
    assign out[2008] = ~(layer_0[129] ^ layer_0[3014]); 
    assign out[2009] = ~(layer_0[453] ^ layer_0[3424]); 
    assign out[2010] = layer_0[3729] ^ layer_0[456]; 
    assign out[2011] = layer_0[2477] ^ layer_0[2263]; 
    assign out[2012] = ~(layer_0[1662] & layer_0[722]); 
    assign out[2013] = layer_0[388] & layer_0[3668]; 
    assign out[2014] = layer_0[2525] | layer_0[3567]; 
    assign out[2015] = ~layer_0[1816]; 
    assign out[2016] = layer_0[2291]; 
    assign out[2017] = ~(layer_0[2620] ^ layer_0[650]); 
    assign out[2018] = ~(layer_0[2578] ^ layer_0[3301]); 
    assign out[2019] = ~(layer_0[1019] ^ layer_0[2571]); 
    assign out[2020] = ~(layer_0[2270] ^ layer_0[2196]); 
    assign out[2021] = layer_0[2482]; 
    assign out[2022] = ~(layer_0[679] | layer_0[1534]); 
    assign out[2023] = layer_0[2504] & ~layer_0[707]; 
    assign out[2024] = ~layer_0[3929] | (layer_0[3929] & layer_0[1017]); 
    assign out[2025] = layer_0[73] & ~layer_0[974]; 
    assign out[2026] = ~(layer_0[2600] ^ layer_0[3738]); 
    assign out[2027] = ~(layer_0[538] ^ layer_0[356]); 
    assign out[2028] = ~layer_0[2238]; 
    assign out[2029] = layer_0[88] & layer_0[3250]; 
    assign out[2030] = layer_0[1735] ^ layer_0[1852]; 
    assign out[2031] = layer_0[2896] & ~layer_0[3630]; 
    assign out[2032] = layer_0[2132] & ~layer_0[622]; 
    assign out[2033] = layer_0[1548]; 
    assign out[2034] = layer_0[3006] ^ layer_0[398]; 
    assign out[2035] = ~(layer_0[3735] & layer_0[187]); 
    assign out[2036] = layer_0[2256] & layer_0[3663]; 
    assign out[2037] = layer_0[863]; 
    assign out[2038] = layer_0[170]; 
    assign out[2039] = layer_0[842] | layer_0[2270]; 
    assign out[2040] = layer_0[1244]; 
    assign out[2041] = ~(layer_0[459] ^ layer_0[2473]); 
    assign out[2042] = ~(layer_0[417] ^ layer_0[2062]); 
    assign out[2043] = ~layer_0[1931] | (layer_0[1931] & layer_0[2421]); 
    assign out[2044] = layer_0[1695] ^ layer_0[2654]; 
    assign out[2045] = ~layer_0[1124]; 
    assign out[2046] = ~(layer_0[2852] ^ layer_0[2757]); 
    assign out[2047] = ~(layer_0[2464] ^ layer_0[469]); 
    assign out[2048] = layer_0[2968] & ~layer_0[3330]; 
    assign out[2049] = layer_0[1944]; 
    assign out[2050] = ~(layer_0[2049] ^ layer_0[316]); 
    assign out[2051] = ~(layer_0[2558] ^ layer_0[1916]); 
    assign out[2052] = ~layer_0[2926]; 
    assign out[2053] = layer_0[2386] ^ layer_0[148]; 
    assign out[2054] = ~layer_0[2334]; 
    assign out[2055] = layer_0[1446] & ~layer_0[3678]; 
    assign out[2056] = layer_0[2509] & ~layer_0[1163]; 
    assign out[2057] = layer_0[1793] ^ layer_0[2054]; 
    assign out[2058] = ~layer_0[3723] | (layer_0[3723] & layer_0[2727]); 
    assign out[2059] = layer_0[520] & ~layer_0[2023]; 
    assign out[2060] = layer_0[1563] ^ layer_0[342]; 
    assign out[2061] = ~(layer_0[2433] | layer_0[920]); 
    assign out[2062] = layer_0[3258] ^ layer_0[3831]; 
    assign out[2063] = layer_0[2283] ^ layer_0[1435]; 
    assign out[2064] = ~(layer_0[220] ^ layer_0[3230]); 
    assign out[2065] = ~layer_0[307]; 
    assign out[2066] = layer_0[1952] ^ layer_0[1183]; 
    assign out[2067] = ~layer_0[605] | (layer_0[347] & layer_0[605]); 
    assign out[2068] = ~(layer_0[3100] ^ layer_0[2535]); 
    assign out[2069] = ~layer_0[1032]; 
    assign out[2070] = ~(layer_0[16] ^ layer_0[326]); 
    assign out[2071] = ~(layer_0[751] ^ layer_0[1507]); 
    assign out[2072] = layer_0[1756] ^ layer_0[212]; 
    assign out[2073] = ~(layer_0[2684] ^ layer_0[2830]); 
    assign out[2074] = layer_0[2041] & ~layer_0[445]; 
    assign out[2075] = layer_0[872] ^ layer_0[3457]; 
    assign out[2076] = ~layer_0[3996]; 
    assign out[2077] = ~layer_0[1337] | (layer_0[1337] & layer_0[1259]); 
    assign out[2078] = layer_0[2678]; 
    assign out[2079] = layer_0[97] ^ layer_0[3821]; 
    assign out[2080] = layer_0[3888] & ~layer_0[1958]; 
    assign out[2081] = layer_0[2262]; 
    assign out[2082] = ~(layer_0[3603] & layer_0[1082]); 
    assign out[2083] = layer_0[3352]; 
    assign out[2084] = layer_0[275]; 
    assign out[2085] = ~(layer_0[2921] & layer_0[3479]); 
    assign out[2086] = ~(layer_0[727] ^ layer_0[1896]); 
    assign out[2087] = layer_0[3419] & layer_0[690]; 
    assign out[2088] = ~(layer_0[855] ^ layer_0[3440]); 
    assign out[2089] = ~(layer_0[3454] | layer_0[1701]); 
    assign out[2090] = layer_0[3307]; 
    assign out[2091] = layer_0[2252] & layer_0[2041]; 
    assign out[2092] = ~layer_0[2656]; 
    assign out[2093] = ~(layer_0[1594] ^ layer_0[481]); 
    assign out[2094] = ~(layer_0[95] | layer_0[1150]); 
    assign out[2095] = layer_0[3544] ^ layer_0[203]; 
    assign out[2096] = layer_0[1895] & layer_0[68]; 
    assign out[2097] = ~(layer_0[289] | layer_0[1904]); 
    assign out[2098] = layer_0[3593] ^ layer_0[1402]; 
    assign out[2099] = layer_0[255] & ~layer_0[960]; 
    assign out[2100] = layer_0[1810] ^ layer_0[3383]; 
    assign out[2101] = layer_0[1639] ^ layer_0[2193]; 
    assign out[2102] = ~(layer_0[1456] ^ layer_0[2986]); 
    assign out[2103] = ~(layer_0[828] ^ layer_0[1626]); 
    assign out[2104] = layer_0[363] ^ layer_0[744]; 
    assign out[2105] = ~(layer_0[3350] ^ layer_0[2622]); 
    assign out[2106] = layer_0[998] ^ layer_0[963]; 
    assign out[2107] = ~layer_0[1125]; 
    assign out[2108] = layer_0[3185] ^ layer_0[1401]; 
    assign out[2109] = layer_0[1889] ^ layer_0[1777]; 
    assign out[2110] = layer_0[3808] ^ layer_0[2035]; 
    assign out[2111] = layer_0[3288] & ~layer_0[3703]; 
    assign out[2112] = layer_0[3444] ^ layer_0[2534]; 
    assign out[2113] = layer_0[1383] & layer_0[3463]; 
    assign out[2114] = layer_0[2160] ^ layer_0[703]; 
    assign out[2115] = layer_0[2347] ^ layer_0[659]; 
    assign out[2116] = ~(layer_0[2798] ^ layer_0[2395]); 
    assign out[2117] = layer_0[157] ^ layer_0[1683]; 
    assign out[2118] = layer_0[1261] ^ layer_0[2289]; 
    assign out[2119] = ~(layer_0[1902] ^ layer_0[2848]); 
    assign out[2120] = ~layer_0[617] | (layer_0[617] & layer_0[2229]); 
    assign out[2121] = ~(layer_0[2798] | layer_0[3448]); 
    assign out[2122] = layer_0[406]; 
    assign out[2123] = layer_0[2634] & ~layer_0[1995]; 
    assign out[2124] = ~layer_0[313] | (layer_0[313] & layer_0[3862]); 
    assign out[2125] = ~(layer_0[422] ^ layer_0[3935]); 
    assign out[2126] = layer_0[3780]; 
    assign out[2127] = layer_0[1348] ^ layer_0[291]; 
    assign out[2128] = ~(layer_0[2117] | layer_0[2923]); 
    assign out[2129] = ~(layer_0[2116] ^ layer_0[574]); 
    assign out[2130] = ~layer_0[1668] | (layer_0[366] & layer_0[1668]); 
    assign out[2131] = ~layer_0[839] | (layer_0[2773] & layer_0[839]); 
    assign out[2132] = ~(layer_0[1092] ^ layer_0[133]); 
    assign out[2133] = ~(layer_0[3261] & layer_0[1016]); 
    assign out[2134] = ~(layer_0[216] & layer_0[1714]); 
    assign out[2135] = ~layer_0[3550]; 
    assign out[2136] = layer_0[1921] ^ layer_0[1722]; 
    assign out[2137] = ~(layer_0[1770] ^ layer_0[3744]); 
    assign out[2138] = ~(layer_0[111] ^ layer_0[2301]); 
    assign out[2139] = layer_0[1993] ^ layer_0[3816]; 
    assign out[2140] = layer_0[485] | layer_0[2907]; 
    assign out[2141] = layer_0[543] ^ layer_0[92]; 
    assign out[2142] = ~(layer_0[932] ^ layer_0[1359]); 
    assign out[2143] = ~layer_0[3655] | (layer_0[3655] & layer_0[1052]); 
    assign out[2144] = layer_0[718]; 
    assign out[2145] = ~layer_0[3456]; 
    assign out[2146] = layer_0[806]; 
    assign out[2147] = layer_0[889]; 
    assign out[2148] = ~(layer_0[1905] ^ layer_0[3705]); 
    assign out[2149] = ~layer_0[579]; 
    assign out[2150] = layer_0[1445]; 
    assign out[2151] = layer_0[3835] ^ layer_0[1718]; 
    assign out[2152] = ~layer_0[2625] | (layer_0[2625] & layer_0[3781]); 
    assign out[2153] = layer_0[1963] & ~layer_0[2596]; 
    assign out[2154] = layer_0[1101] & layer_0[2219]; 
    assign out[2155] = ~(layer_0[3805] ^ layer_0[3814]); 
    assign out[2156] = layer_0[318]; 
    assign out[2157] = layer_0[3382]; 
    assign out[2158] = ~(layer_0[3687] ^ layer_0[1799]); 
    assign out[2159] = layer_0[403] ^ layer_0[3681]; 
    assign out[2160] = ~layer_0[833]; 
    assign out[2161] = layer_0[1375] & ~layer_0[1462]; 
    assign out[2162] = layer_0[2721] ^ layer_0[1851]; 
    assign out[2163] = ~(layer_0[950] ^ layer_0[2734]); 
    assign out[2164] = layer_0[3007] ^ layer_0[3859]; 
    assign out[2165] = layer_0[3529] | layer_0[2084]; 
    assign out[2166] = ~(layer_0[2428] ^ layer_0[2063]); 
    assign out[2167] = layer_0[2366] ^ layer_0[3829]; 
    assign out[2168] = ~(layer_0[3907] ^ layer_0[3142]); 
    assign out[2169] = layer_0[82]; 
    assign out[2170] = ~layer_0[164]; 
    assign out[2171] = layer_0[1614] & layer_0[2271]; 
    assign out[2172] = ~layer_0[2689]; 
    assign out[2173] = layer_0[3326] ^ layer_0[3337]; 
    assign out[2174] = ~layer_0[1307] | (layer_0[1307] & layer_0[3303]); 
    assign out[2175] = layer_0[1817] ^ layer_0[3370]; 
    assign out[2176] = ~(layer_0[3051] ^ layer_0[1769]); 
    assign out[2177] = ~(layer_0[2021] ^ layer_0[1542]); 
    assign out[2178] = layer_0[2588] & ~layer_0[2221]; 
    assign out[2179] = ~layer_0[2327]; 
    assign out[2180] = ~layer_0[902] | (layer_0[902] & layer_0[3195]); 
    assign out[2181] = layer_0[667]; 
    assign out[2182] = layer_0[343] & ~layer_0[2203]; 
    assign out[2183] = ~(layer_0[3813] ^ layer_0[886]); 
    assign out[2184] = ~(layer_0[1434] ^ layer_0[1394]); 
    assign out[2185] = layer_0[854] & layer_0[1167]; 
    assign out[2186] = ~(layer_0[2833] ^ layer_0[2190]); 
    assign out[2187] = ~layer_0[2667] | (layer_0[2417] & layer_0[2667]); 
    assign out[2188] = ~(layer_0[2853] | layer_0[530]); 
    assign out[2189] = layer_0[3136] | layer_0[2471]; 
    assign out[2190] = layer_0[2243] | layer_0[3059]; 
    assign out[2191] = ~layer_0[629] | (layer_0[2408] & layer_0[629]); 
    assign out[2192] = ~(layer_0[265] & layer_0[3067]); 
    assign out[2193] = layer_0[206] ^ layer_0[591]; 
    assign out[2194] = ~(layer_0[3104] ^ layer_0[1299]); 
    assign out[2195] = ~layer_0[1378] | (layer_0[1378] & layer_0[2516]); 
    assign out[2196] = ~(layer_0[968] ^ layer_0[1679]); 
    assign out[2197] = layer_0[1222] | layer_0[2985]; 
    assign out[2198] = layer_0[3132] ^ layer_0[2822]; 
    assign out[2199] = ~(layer_0[1552] ^ layer_0[3833]); 
    assign out[2200] = layer_0[1392] ^ layer_0[479]; 
    assign out[2201] = ~layer_0[578]; 
    assign out[2202] = ~(layer_0[3449] | layer_0[1676]); 
    assign out[2203] = layer_0[446] & ~layer_0[694]; 
    assign out[2204] = layer_0[3855] & layer_0[2951]; 
    assign out[2205] = layer_0[715] ^ layer_0[2792]; 
    assign out[2206] = layer_0[2829] ^ layer_0[3078]; 
    assign out[2207] = ~(layer_0[3616] ^ layer_0[1067]); 
    assign out[2208] = layer_0[1949] | layer_0[326]; 
    assign out[2209] = layer_0[2090] ^ layer_0[2]; 
    assign out[2210] = layer_0[2025] ^ layer_0[2312]; 
    assign out[2211] = ~layer_0[1900] | (layer_0[160] & layer_0[1900]); 
    assign out[2212] = ~layer_0[918] | (layer_0[918] & layer_0[3806]); 
    assign out[2213] = ~layer_0[189]; 
    assign out[2214] = ~layer_0[44] | (layer_0[2155] & layer_0[44]); 
    assign out[2215] = ~(layer_0[2930] ^ layer_0[691]); 
    assign out[2216] = ~(layer_0[3495] ^ layer_0[632]); 
    assign out[2217] = ~(layer_0[1213] ^ layer_0[1449]); 
    assign out[2218] = ~(layer_0[3793] ^ layer_0[555]); 
    assign out[2219] = ~(layer_0[800] ^ layer_0[3166]); 
    assign out[2220] = layer_0[1494]; 
    assign out[2221] = layer_0[3126]; 
    assign out[2222] = ~layer_0[3012]; 
    assign out[2223] = layer_0[185] ^ layer_0[433]; 
    assign out[2224] = layer_0[3341] ^ layer_0[1258]; 
    assign out[2225] = layer_0[731] ^ layer_0[1431]; 
    assign out[2226] = layer_0[812] & layer_0[709]; 
    assign out[2227] = layer_0[154] ^ layer_0[2714]; 
    assign out[2228] = ~(layer_0[3129] ^ layer_0[603]); 
    assign out[2229] = layer_0[1864] ^ layer_0[1796]; 
    assign out[2230] = ~(layer_0[1663] ^ layer_0[1600]); 
    assign out[2231] = ~layer_0[569]; 
    assign out[2232] = layer_0[1459] ^ layer_0[3079]; 
    assign out[2233] = layer_0[283]; 
    assign out[2234] = layer_0[3420]; 
    assign out[2235] = ~(layer_0[1774] ^ layer_0[381]); 
    assign out[2236] = ~(layer_0[3131] ^ layer_0[3860]); 
    assign out[2237] = layer_0[425] & layer_0[624]; 
    assign out[2238] = ~(layer_0[3900] ^ layer_0[3015]); 
    assign out[2239] = ~layer_0[2363] | (layer_0[3596] & layer_0[2363]); 
    assign out[2240] = layer_0[2338] ^ layer_0[2425]; 
    assign out[2241] = ~layer_0[3552] | (layer_0[3552] & layer_0[204]); 
    assign out[2242] = ~layer_0[277]; 
    assign out[2243] = layer_0[2606] ^ layer_0[2808]; 
    assign out[2244] = ~(layer_0[1726] | layer_0[3449]); 
    assign out[2245] = layer_0[1663] ^ layer_0[2916]; 
    assign out[2246] = ~layer_0[2104]; 
    assign out[2247] = ~(layer_0[2631] ^ layer_0[2174]); 
    assign out[2248] = ~layer_0[1480]; 
    assign out[2249] = ~(layer_0[1943] | layer_0[2022]); 
    assign out[2250] = ~(layer_0[1001] ^ layer_0[3754]); 
    assign out[2251] = ~layer_0[2055]; 
    assign out[2252] = layer_0[3075] & ~layer_0[2414]; 
    assign out[2253] = layer_0[3200]; 
    assign out[2254] = ~(layer_0[2396] | layer_0[1965]); 
    assign out[2255] = ~(layer_0[3386] ^ layer_0[2702]); 
    assign out[2256] = ~layer_0[3532] | (layer_0[12] & layer_0[3532]); 
    assign out[2257] = layer_0[1599] | layer_0[1498]; 
    assign out[2258] = layer_0[1175]; 
    assign out[2259] = layer_0[2800] ^ layer_0[3418]; 
    assign out[2260] = layer_0[3507] ^ layer_0[3614]; 
    assign out[2261] = ~layer_0[466] | (layer_0[510] & layer_0[466]); 
    assign out[2262] = ~layer_0[3022]; 
    assign out[2263] = ~layer_0[3074]; 
    assign out[2264] = layer_0[756] ^ layer_0[2289]; 
    assign out[2265] = layer_0[2780]; 
    assign out[2266] = ~(layer_0[3548] & layer_0[2012]); 
    assign out[2267] = layer_0[29]; 
    assign out[2268] = ~(layer_0[1873] ^ layer_0[3438]); 
    assign out[2269] = layer_0[3477]; 
    assign out[2270] = layer_0[2047] & ~layer_0[2953]; 
    assign out[2271] = ~(layer_0[1807] ^ layer_0[2517]); 
    assign out[2272] = layer_0[915] ^ layer_0[1961]; 
    assign out[2273] = layer_0[280] ^ layer_0[2284]; 
    assign out[2274] = ~(layer_0[1549] ^ layer_0[3643]); 
    assign out[2275] = layer_0[115] ^ layer_0[2179]; 
    assign out[2276] = layer_0[851] ^ layer_0[845]; 
    assign out[2277] = ~layer_0[577]; 
    assign out[2278] = layer_0[475]; 
    assign out[2279] = ~(layer_0[3774] ^ layer_0[1857]); 
    assign out[2280] = ~layer_0[2336]; 
    assign out[2281] = layer_0[2642] & layer_0[2932]; 
    assign out[2282] = ~(layer_0[1100] ^ layer_0[2908]); 
    assign out[2283] = layer_0[2232] ^ layer_0[1350]; 
    assign out[2284] = ~(layer_0[584] ^ layer_0[2991]); 
    assign out[2285] = ~layer_0[947]; 
    assign out[2286] = layer_0[2906]; 
    assign out[2287] = ~(layer_0[3050] | layer_0[650]); 
    assign out[2288] = layer_0[2825] ^ layer_0[2492]; 
    assign out[2289] = ~(layer_0[3367] ^ layer_0[1322]); 
    assign out[2290] = ~(layer_0[1302] ^ layer_0[237]); 
    assign out[2291] = ~(layer_0[79] ^ layer_0[1898]); 
    assign out[2292] = layer_0[43]; 
    assign out[2293] = layer_0[2404] ^ layer_0[3748]; 
    assign out[2294] = layer_0[721] ^ layer_0[3605]; 
    assign out[2295] = layer_0[195] & layer_0[2217]; 
    assign out[2296] = layer_0[1328] ^ layer_0[1115]; 
    assign out[2297] = layer_0[2781]; 
    assign out[2298] = ~(layer_0[3618] ^ layer_0[1803]); 
    assign out[2299] = layer_0[370] & layer_0[2694]; 
    assign out[2300] = layer_0[1280]; 
    assign out[2301] = ~layer_0[1455]; 
    assign out[2302] = layer_0[1536] ^ layer_0[2375]; 
    assign out[2303] = layer_0[382] & ~layer_0[3153]; 
    assign out[2304] = layer_0[2423] ^ layer_0[1818]; 
    assign out[2305] = layer_0[3220] ^ layer_0[3615]; 
    assign out[2306] = ~(layer_0[1186] ^ layer_0[3455]); 
    assign out[2307] = layer_0[3800] & layer_0[2109]; 
    assign out[2308] = layer_0[2563] ^ layer_0[3989]; 
    assign out[2309] = layer_0[1300] ^ layer_0[1677]; 
    assign out[2310] = layer_0[484] ^ layer_0[358]; 
    assign out[2311] = ~(layer_0[944] ^ layer_0[174]); 
    assign out[2312] = layer_0[970] ^ layer_0[887]; 
    assign out[2313] = ~(layer_0[1492] | layer_0[244]); 
    assign out[2314] = layer_0[1209] & ~layer_0[1772]; 
    assign out[2315] = ~layer_0[2593]; 
    assign out[2316] = layer_0[1154]; 
    assign out[2317] = ~(layer_0[2493] ^ layer_0[369]); 
    assign out[2318] = ~(layer_0[123] & layer_0[3265]); 
    assign out[2319] = ~(layer_0[3803] ^ layer_0[1032]); 
    assign out[2320] = ~(layer_0[2782] ^ layer_0[424]); 
    assign out[2321] = layer_0[463] & ~layer_0[1717]; 
    assign out[2322] = layer_0[2146] ^ layer_0[3031]; 
    assign out[2323] = ~(layer_0[2232] & layer_0[1598]); 
    assign out[2324] = ~(layer_0[2409] ^ layer_0[3101]); 
    assign out[2325] = layer_0[1264] & layer_0[506]; 
    assign out[2326] = layer_0[2141] & ~layer_0[720]; 
    assign out[2327] = layer_0[3511] ^ layer_0[2359]; 
    assign out[2328] = layer_0[131] & layer_0[797]; 
    assign out[2329] = layer_0[3048] & layer_0[3228]; 
    assign out[2330] = layer_0[2748] ^ layer_0[1504]; 
    assign out[2331] = layer_0[643] & ~layer_0[1846]; 
    assign out[2332] = layer_0[3530] ^ layer_0[2149]; 
    assign out[2333] = ~layer_0[334]; 
    assign out[2334] = layer_0[2730] & layer_0[2302]; 
    assign out[2335] = ~layer_0[540]; 
    assign out[2336] = ~(layer_0[3747] ^ layer_0[1759]); 
    assign out[2337] = ~layer_0[1253] | (layer_0[2739] & layer_0[1253]); 
    assign out[2338] = layer_0[2863] & layer_0[3894]; 
    assign out[2339] = ~(layer_0[1325] | layer_0[3329]); 
    assign out[2340] = ~(layer_0[3306] ^ layer_0[400]); 
    assign out[2341] = ~(layer_0[3864] | layer_0[3971]); 
    assign out[2342] = ~(layer_0[3591] | layer_0[251]); 
    assign out[2343] = layer_0[1073] ^ layer_0[67]; 
    assign out[2344] = layer_0[2300]; 
    assign out[2345] = ~layer_0[2575]; 
    assign out[2346] = ~(layer_0[3123] ^ layer_0[387]); 
    assign out[2347] = layer_0[3564] | layer_0[1102]; 
    assign out[2348] = ~layer_0[2575]; 
    assign out[2349] = ~(layer_0[1928] ^ layer_0[1664]); 
    assign out[2350] = layer_0[3562] & ~layer_0[2646]; 
    assign out[2351] = ~(layer_0[2153] ^ layer_0[1004]); 
    assign out[2352] = layer_0[2545]; 
    assign out[2353] = ~(layer_0[774] ^ layer_0[3079]); 
    assign out[2354] = layer_0[3922] & layer_0[1820]; 
    assign out[2355] = layer_0[176] ^ layer_0[3473]; 
    assign out[2356] = ~(layer_0[1470] ^ layer_0[1013]); 
    assign out[2357] = ~layer_0[2206]; 
    assign out[2358] = ~layer_0[3375]; 
    assign out[2359] = ~layer_0[675] | (layer_0[675] & layer_0[2738]); 
    assign out[2360] = ~(layer_0[3767] ^ layer_0[2048]); 
    assign out[2361] = layer_0[912]; 
    assign out[2362] = ~(layer_0[1863] ^ layer_0[1547]); 
    assign out[2363] = layer_0[2371] & ~layer_0[2976]; 
    assign out[2364] = ~layer_0[2875] | (layer_0[2875] & layer_0[3106]); 
    assign out[2365] = layer_0[1288]; 
    assign out[2366] = ~(layer_0[3047] ^ layer_0[2540]); 
    assign out[2367] = ~(layer_0[3884] ^ layer_0[715]); 
    assign out[2368] = layer_0[3032] ^ layer_0[1777]; 
    assign out[2369] = ~layer_0[2769] | (layer_0[3321] & layer_0[2769]); 
    assign out[2370] = ~(layer_0[394] ^ layer_0[1858]); 
    assign out[2371] = layer_0[858] & layer_0[2544]; 
    assign out[2372] = layer_0[2444] ^ layer_0[1892]; 
    assign out[2373] = ~(layer_0[130] ^ layer_0[637]); 
    assign out[2374] = layer_0[3930] & ~layer_0[2057]; 
    assign out[2375] = ~(layer_0[3121] ^ layer_0[3972]); 
    assign out[2376] = layer_0[2607] & ~layer_0[1597]; 
    assign out[2377] = ~layer_0[350]; 
    assign out[2378] = ~layer_0[2663]; 
    assign out[2379] = ~layer_0[1128]; 
    assign out[2380] = ~(layer_0[1474] ^ layer_0[3736]); 
    assign out[2381] = layer_0[1790]; 
    assign out[2382] = layer_0[2461] & ~layer_0[1109]; 
    assign out[2383] = ~(layer_0[1120] ^ layer_0[1287]); 
    assign out[2384] = ~layer_0[3450]; 
    assign out[2385] = ~(layer_0[3369] ^ layer_0[136]); 
    assign out[2386] = ~(layer_0[3471] ^ layer_0[1826]); 
    assign out[2387] = layer_0[113] ^ layer_0[1750]; 
    assign out[2388] = layer_0[83] ^ layer_0[472]; 
    assign out[2389] = layer_0[3873]; 
    assign out[2390] = ~layer_0[2985]; 
    assign out[2391] = layer_0[201]; 
    assign out[2392] = ~(layer_0[729] | layer_0[1727]); 
    assign out[2393] = layer_0[3924] ^ layer_0[1878]; 
    assign out[2394] = layer_0[3110] & ~layer_0[1772]; 
    assign out[2395] = layer_0[3446] ^ layer_0[1447]; 
    assign out[2396] = layer_0[3585] & ~layer_0[1570]; 
    assign out[2397] = layer_0[3988] & layer_0[3954]; 
    assign out[2398] = layer_0[2955] ^ layer_0[2031]; 
    assign out[2399] = layer_0[801] ^ layer_0[770]; 
    assign out[2400] = layer_0[2345] ^ layer_0[3085]; 
    assign out[2401] = layer_0[3998]; 
    assign out[2402] = layer_0[1747]; 
    assign out[2403] = layer_0[1403] & layer_0[2056]; 
    assign out[2404] = layer_0[1371] & ~layer_0[3990]; 
    assign out[2405] = ~(layer_0[1637] ^ layer_0[2620]); 
    assign out[2406] = ~layer_0[1170]; 
    assign out[2407] = layer_0[699] & layer_0[2635]; 
    assign out[2408] = layer_0[3289] ^ layer_0[3235]; 
    assign out[2409] = ~(layer_0[1546] ^ layer_0[2501]); 
    assign out[2410] = ~(layer_0[1665] ^ layer_0[2886]); 
    assign out[2411] = ~(layer_0[1823] ^ layer_0[74]); 
    assign out[2412] = layer_0[2918] ^ layer_0[2283]; 
    assign out[2413] = ~(layer_0[2259] ^ layer_0[747]); 
    assign out[2414] = layer_0[869]; 
    assign out[2415] = ~(layer_0[1196] | layer_0[3965]); 
    assign out[2416] = layer_0[2186] ^ layer_0[1613]; 
    assign out[2417] = layer_0[1571] ^ layer_0[752]; 
    assign out[2418] = ~(layer_0[2947] ^ layer_0[3744]); 
    assign out[2419] = ~(layer_0[3035] | layer_0[3197]); 
    assign out[2420] = layer_0[69] ^ layer_0[2621]; 
    assign out[2421] = layer_0[905] ^ layer_0[848]; 
    assign out[2422] = ~(layer_0[3853] | layer_0[1540]); 
    assign out[2423] = ~(layer_0[1923] ^ layer_0[3055]); 
    assign out[2424] = ~layer_0[791] | (layer_0[791] & layer_0[1956]); 
    assign out[2425] = ~(layer_0[1292] | layer_0[2619]); 
    assign out[2426] = layer_0[2435] & ~layer_0[1420]; 
    assign out[2427] = layer_0[3818] ^ layer_0[3348]; 
    assign out[2428] = layer_0[1189] ^ layer_0[2806]; 
    assign out[2429] = layer_0[2368] & ~layer_0[3909]; 
    assign out[2430] = layer_0[2488]; 
    assign out[2431] = ~layer_0[3138]; 
    assign out[2432] = layer_0[1464]; 
    assign out[2433] = layer_0[3398] ^ layer_0[1424]; 
    assign out[2434] = ~layer_0[1888]; 
    assign out[2435] = layer_0[3837]; 
    assign out[2436] = ~(layer_0[2831] ^ layer_0[1860]); 
    assign out[2437] = ~layer_0[1188]; 
    assign out[2438] = layer_0[2613] ^ layer_0[3751]; 
    assign out[2439] = ~(layer_0[1264] ^ layer_0[716]); 
    assign out[2440] = ~(layer_0[734] ^ layer_0[161]); 
    assign out[2441] = ~(layer_0[1608] ^ layer_0[3285]); 
    assign out[2442] = layer_0[3216]; 
    assign out[2443] = ~layer_0[1094]; 
    assign out[2444] = ~layer_0[477]; 
    assign out[2445] = layer_0[3088] ^ layer_0[1456]; 
    assign out[2446] = layer_0[3953] ^ layer_0[339]; 
    assign out[2447] = layer_0[3727] ^ layer_0[1192]; 
    assign out[2448] = ~(layer_0[2425] | layer_0[2015]); 
    assign out[2449] = layer_0[151] ^ layer_0[2742]; 
    assign out[2450] = ~(layer_0[276] ^ layer_0[3034]); 
    assign out[2451] = layer_0[1241] ^ layer_0[71]; 
    assign out[2452] = layer_0[1062] ^ layer_0[1655]; 
    assign out[2453] = layer_0[1588]; 
    assign out[2454] = layer_0[2169] ^ layer_0[1981]; 
    assign out[2455] = ~layer_0[2269]; 
    assign out[2456] = ~layer_0[103] | (layer_0[2519] & layer_0[103]); 
    assign out[2457] = ~layer_0[1479]; 
    assign out[2458] = ~(layer_0[1180] ^ layer_0[2822]); 
    assign out[2459] = layer_0[2611] & ~layer_0[354]; 
    assign out[2460] = layer_0[78] & ~layer_0[215]; 
    assign out[2461] = layer_0[3549] ^ layer_0[573]; 
    assign out[2462] = layer_0[264] & ~layer_0[3499]; 
    assign out[2463] = layer_0[2962] & ~layer_0[3001]; 
    assign out[2464] = layer_0[3957] ^ layer_0[63]; 
    assign out[2465] = layer_0[1826] ^ layer_0[2595]; 
    assign out[2466] = layer_0[3095] & layer_0[2740]; 
    assign out[2467] = ~(layer_0[348] ^ layer_0[2917]); 
    assign out[2468] = layer_0[2877] & ~layer_0[1214]; 
    assign out[2469] = layer_0[2473] & layer_0[784]; 
    assign out[2470] = ~layer_0[3261]; 
    assign out[2471] = layer_0[2877] & ~layer_0[3189]; 
    assign out[2472] = ~layer_0[5]; 
    assign out[2473] = ~(layer_0[495] | layer_0[2587]); 
    assign out[2474] = ~layer_0[3057]; 
    assign out[2475] = ~(layer_0[3963] ^ layer_0[1635]); 
    assign out[2476] = layer_0[908] ^ layer_0[994]; 
    assign out[2477] = layer_0[1647] ^ layer_0[3869]; 
    assign out[2478] = layer_0[2922] & ~layer_0[1929]; 
    assign out[2479] = layer_0[3828] ^ layer_0[1913]; 
    assign out[2480] = ~layer_0[698]; 
    assign out[2481] = layer_0[2796]; 
    assign out[2482] = ~(layer_0[3429] ^ layer_0[2165]); 
    assign out[2483] = ~(layer_0[3944] ^ layer_0[1742]); 
    assign out[2484] = ~(layer_0[3199] ^ layer_0[3204]); 
    assign out[2485] = ~(layer_0[575] ^ layer_0[911]); 
    assign out[2486] = ~layer_0[3253]; 
    assign out[2487] = layer_0[2959] | layer_0[2965]; 
    assign out[2488] = layer_0[1185] ^ layer_0[2574]; 
    assign out[2489] = ~layer_0[1478]; 
    assign out[2490] = layer_0[3492]; 
    assign out[2491] = ~(layer_0[1873] ^ layer_0[647]); 
    assign out[2492] = ~(layer_0[1645] ^ layer_0[118]); 
    assign out[2493] = layer_0[2174]; 
    assign out[2494] = ~(layer_0[3361] | layer_0[1396]); 
    assign out[2495] = ~(layer_0[2224] ^ layer_0[2488]); 
    assign out[2496] = layer_0[1585] & ~layer_0[2194]; 
    assign out[2497] = layer_0[3373] & layer_0[2348]; 
    assign out[2498] = layer_0[2085]; 
    assign out[2499] = layer_0[3658] & layer_0[946]; 
    assign out[2500] = ~(layer_0[3422] ^ layer_0[2009]); 
    assign out[2501] = layer_0[3903] & ~layer_0[184]; 
    assign out[2502] = layer_0[1704] & layer_0[826]; 
    assign out[2503] = layer_0[760] ^ layer_0[2851]; 
    assign out[2504] = layer_0[2668] & ~layer_0[974]; 
    assign out[2505] = layer_0[3734] & ~layer_0[31]; 
    assign out[2506] = ~layer_0[2430] | (layer_0[2724] & layer_0[2430]); 
    assign out[2507] = layer_0[2046] & ~layer_0[1066]; 
    assign out[2508] = ~layer_0[3648]; 
    assign out[2509] = layer_0[2214] ^ layer_0[2760]; 
    assign out[2510] = ~layer_0[2290]; 
    assign out[2511] = layer_0[1018] ^ layer_0[3865]; 
    assign out[2512] = ~(layer_0[540] ^ layer_0[2772]); 
    assign out[2513] = ~(layer_0[745] ^ layer_0[2824]); 
    assign out[2514] = ~(layer_0[3619] ^ layer_0[3563]); 
    assign out[2515] = layer_0[3260]; 
    assign out[2516] = layer_0[461]; 
    assign out[2517] = layer_0[3390] ^ layer_0[2859]; 
    assign out[2518] = layer_0[1586]; 
    assign out[2519] = ~layer_0[378] | (layer_0[378] & layer_0[3356]); 
    assign out[2520] = layer_0[3382]; 
    assign out[2521] = ~layer_0[2343]; 
    assign out[2522] = layer_0[1335] ^ layer_0[1357]; 
    assign out[2523] = layer_0[1193] | layer_0[3801]; 
    assign out[2524] = layer_0[3016] | layer_0[2173]; 
    assign out[2525] = ~(layer_0[1004] ^ layer_0[1765]); 
    assign out[2526] = ~(layer_0[1040] ^ layer_0[3923]); 
    assign out[2527] = layer_0[3241] & layer_0[1349]; 
    assign out[2528] = ~(layer_0[1079] ^ layer_0[3214]); 
    assign out[2529] = layer_0[3759]; 
    assign out[2530] = layer_0[329] ^ layer_0[712]; 
    assign out[2531] = ~(layer_0[3715] ^ layer_0[933]); 
    assign out[2532] = ~(layer_0[2195] ^ layer_0[888]); 
    assign out[2533] = layer_0[804]; 
    assign out[2534] = layer_0[1854] ^ layer_0[693]; 
    assign out[2535] = ~(layer_0[1607] ^ layer_0[1372]); 
    assign out[2536] = ~(layer_0[3526] & layer_0[3317]); 
    assign out[2537] = layer_0[894] ^ layer_0[2076]; 
    assign out[2538] = layer_0[966] ^ layer_0[1244]; 
    assign out[2539] = layer_0[3659]; 
    assign out[2540] = ~layer_0[3155] | (layer_0[3155] & layer_0[1509]); 
    assign out[2541] = layer_0[3165] & ~layer_0[2638]; 
    assign out[2542] = ~(layer_0[128] & layer_0[2392]); 
    assign out[2543] = layer_0[3625] | layer_0[2633]; 
    assign out[2544] = layer_0[58] & ~layer_0[2716]; 
    assign out[2545] = layer_0[2052] & ~layer_0[2638]; 
    assign out[2546] = ~layer_0[3525]; 
    assign out[2547] = layer_0[3674]; 
    assign out[2548] = ~(layer_0[3232] ^ layer_0[533]); 
    assign out[2549] = layer_0[1634]; 
    assign out[2550] = 1'b0; 
    assign out[2551] = 1'b0; 
    assign out[2552] = 1'b0; 
    assign out[2553] = 1'b0; 
    assign out[2554] = 1'b0; 
    assign out[2555] = 1'b0; 
    assign out[2556] = 1'b0; 
    assign out[2557] = 1'b0; 
    assign out[2558] = 1'b0; 
    assign out[2559] = 1'b0; 
    assign out[2560] = 1'b0; 
    assign out[2561] = 1'b0; 
    assign out[2562] = 1'b0; 
    assign out[2563] = 1'b0; 
    assign out[2564] = 1'b0; 
    assign out[2565] = 1'b0; 
    assign out[2566] = 1'b0; 
    assign out[2567] = 1'b0; 
    assign out[2568] = 1'b0; 
    assign out[2569] = 1'b0; 
    assign out[2570] = 1'b0; 
    assign out[2571] = 1'b0; 
    assign out[2572] = 1'b0; 
    assign out[2573] = 1'b0; 
    assign out[2574] = 1'b0; 
    assign out[2575] = 1'b0; 
    assign out[2576] = 1'b0; 
    assign out[2577] = 1'b0; 
    assign out[2578] = 1'b0; 
    assign out[2579] = 1'b0; 
    assign out[2580] = 1'b0; 
    assign out[2581] = 1'b0; 
    assign out[2582] = 1'b0; 
    assign out[2583] = 1'b0; 
    assign out[2584] = 1'b0; 
    assign out[2585] = 1'b0; 
    assign out[2586] = 1'b0; 
    assign out[2587] = 1'b0; 
    assign out[2588] = 1'b0; 
    assign out[2589] = 1'b0; 
    assign out[2590] = 1'b0; 
    assign out[2591] = 1'b0; 
    assign out[2592] = 1'b0; 
    assign out[2593] = 1'b0; 
    assign out[2594] = 1'b0; 
    assign out[2595] = 1'b0; 
    assign out[2596] = 1'b0; 
    assign out[2597] = 1'b0; 
    assign out[2598] = 1'b0; 
    assign out[2599] = 1'b0; 
    assign out[2600] = 1'b0; 
    assign out[2601] = 1'b0; 
    assign out[2602] = 1'b0; 
    assign out[2603] = 1'b0; 
    assign out[2604] = 1'b0; 
    assign out[2605] = 1'b0; 
    assign out[2606] = 1'b0; 
    assign out[2607] = 1'b0; 
    assign out[2608] = 1'b0; 
    assign out[2609] = 1'b0; 
    assign out[2610] = 1'b0; 
    assign out[2611] = 1'b0; 
    assign out[2612] = 1'b0; 
    assign out[2613] = 1'b0; 
    assign out[2614] = 1'b0; 
    assign out[2615] = 1'b0; 
    assign out[2616] = 1'b0; 
    assign out[2617] = 1'b0; 
    assign out[2618] = 1'b0; 
    assign out[2619] = 1'b0; 
    assign out[2620] = 1'b0; 
    assign out[2621] = 1'b0; 
    assign out[2622] = 1'b0; 
    assign out[2623] = 1'b0; 
    assign out[2624] = 1'b0; 
    assign out[2625] = 1'b0; 
    assign out[2626] = 1'b0; 
    assign out[2627] = 1'b0; 
    assign out[2628] = 1'b0; 
    assign out[2629] = 1'b0; 
    assign out[2630] = 1'b0; 
    assign out[2631] = 1'b0; 
    assign out[2632] = 1'b0; 
    assign out[2633] = 1'b0; 
    assign out[2634] = 1'b0; 
    assign out[2635] = 1'b0; 
    assign out[2636] = 1'b0; 
    assign out[2637] = 1'b0; 
    assign out[2638] = 1'b0; 
    assign out[2639] = 1'b0; 
    assign out[2640] = 1'b0; 
    assign out[2641] = 1'b0; 
    assign out[2642] = 1'b0; 
    assign out[2643] = 1'b0; 
    assign out[2644] = 1'b0; 
    assign out[2645] = 1'b0; 
    assign out[2646] = 1'b0; 
    assign out[2647] = 1'b0; 
    assign out[2648] = 1'b0; 
    assign out[2649] = 1'b0; 
    assign out[2650] = 1'b0; 
    assign out[2651] = 1'b0; 
    assign out[2652] = 1'b0; 
    assign out[2653] = 1'b0; 
    assign out[2654] = 1'b0; 
    assign out[2655] = 1'b0; 
    assign out[2656] = 1'b0; 
    assign out[2657] = 1'b0; 
    assign out[2658] = 1'b0; 
    assign out[2659] = 1'b0; 
    assign out[2660] = 1'b0; 
    assign out[2661] = 1'b0; 
    assign out[2662] = 1'b0; 
    assign out[2663] = 1'b0; 
    assign out[2664] = 1'b0; 
    assign out[2665] = 1'b0; 
    assign out[2666] = 1'b0; 
    assign out[2667] = 1'b0; 
    assign out[2668] = 1'b0; 
    assign out[2669] = 1'b0; 
    assign out[2670] = 1'b0; 
    assign out[2671] = 1'b0; 
    assign out[2672] = 1'b0; 
    assign out[2673] = 1'b0; 
    assign out[2674] = 1'b0; 
    assign out[2675] = 1'b0; 
    assign out[2676] = 1'b0; 
    assign out[2677] = 1'b0; 
    assign out[2678] = 1'b0; 
    assign out[2679] = 1'b0; 
    assign out[2680] = 1'b0; 
    assign out[2681] = 1'b0; 
    assign out[2682] = 1'b0; 
    assign out[2683] = 1'b0; 
    assign out[2684] = 1'b0; 
    assign out[2685] = 1'b0; 
    assign out[2686] = 1'b0; 
    assign out[2687] = 1'b0; 
    assign out[2688] = 1'b0; 
    assign out[2689] = 1'b0; 
    assign out[2690] = 1'b0; 
    assign out[2691] = 1'b0; 
    assign out[2692] = 1'b0; 
    assign out[2693] = 1'b0; 
    assign out[2694] = 1'b0; 
    assign out[2695] = 1'b0; 
    assign out[2696] = 1'b0; 
    assign out[2697] = 1'b0; 
    assign out[2698] = 1'b0; 
    assign out[2699] = 1'b0; 
    assign out[2700] = 1'b0; 
    assign out[2701] = 1'b0; 
    assign out[2702] = 1'b0; 
    assign out[2703] = 1'b0; 
    assign out[2704] = 1'b0; 
    assign out[2705] = 1'b0; 
    assign out[2706] = 1'b0; 
    assign out[2707] = 1'b0; 
    assign out[2708] = 1'b0; 
    assign out[2709] = 1'b0; 
    assign out[2710] = 1'b0; 
    assign out[2711] = 1'b0; 
    assign out[2712] = 1'b0; 
    assign out[2713] = 1'b0; 
    assign out[2714] = 1'b0; 
    assign out[2715] = 1'b0; 
    assign out[2716] = 1'b0; 
    assign out[2717] = 1'b0; 
    assign out[2718] = 1'b0; 
    assign out[2719] = 1'b0; 
    assign out[2720] = 1'b0; 
    assign out[2721] = 1'b0; 
    assign out[2722] = 1'b0; 
    assign out[2723] = 1'b0; 
    assign out[2724] = 1'b0; 
    assign out[2725] = 1'b0; 
    assign out[2726] = 1'b0; 
    assign out[2727] = 1'b0; 
    assign out[2728] = 1'b0; 
    assign out[2729] = 1'b0; 
    assign out[2730] = 1'b0; 
    assign out[2731] = 1'b0; 
    assign out[2732] = 1'b0; 
    assign out[2733] = 1'b0; 
    assign out[2734] = 1'b0; 
    assign out[2735] = 1'b0; 
    assign out[2736] = 1'b0; 
    assign out[2737] = 1'b0; 
    assign out[2738] = 1'b0; 
    assign out[2739] = 1'b0; 
    assign out[2740] = 1'b0; 
    assign out[2741] = 1'b0; 
    assign out[2742] = 1'b0; 
    assign out[2743] = 1'b0; 
    assign out[2744] = 1'b0; 
    assign out[2745] = 1'b0; 
    assign out[2746] = 1'b0; 
    assign out[2747] = 1'b0; 
    assign out[2748] = 1'b0; 
    assign out[2749] = 1'b0; 
    assign out[2750] = 1'b0; 
    assign out[2751] = 1'b0; 
    assign out[2752] = 1'b0; 
    assign out[2753] = 1'b0; 
    assign out[2754] = 1'b0; 
    assign out[2755] = 1'b0; 
    assign out[2756] = 1'b0; 
    assign out[2757] = 1'b0; 
    assign out[2758] = 1'b0; 
    assign out[2759] = 1'b0; 
    assign out[2760] = 1'b0; 
    assign out[2761] = 1'b0; 
    assign out[2762] = 1'b0; 
    assign out[2763] = 1'b0; 
    assign out[2764] = 1'b0; 
    assign out[2765] = 1'b0; 
    assign out[2766] = 1'b0; 
    assign out[2767] = 1'b0; 
    assign out[2768] = 1'b0; 
    assign out[2769] = 1'b0; 
    assign out[2770] = 1'b0; 
    assign out[2771] = 1'b0; 
    assign out[2772] = 1'b0; 
    assign out[2773] = 1'b0; 
    assign out[2774] = 1'b0; 
    assign out[2775] = 1'b0; 
    assign out[2776] = 1'b0; 
    assign out[2777] = 1'b0; 
    assign out[2778] = 1'b0; 
    assign out[2779] = 1'b0; 
    assign out[2780] = 1'b0; 
    assign out[2781] = 1'b0; 
    assign out[2782] = 1'b0; 
    assign out[2783] = 1'b0; 
    assign out[2784] = 1'b0; 
    assign out[2785] = 1'b0; 
    assign out[2786] = 1'b0; 
    assign out[2787] = 1'b0; 
    assign out[2788] = 1'b0; 
    assign out[2789] = 1'b0; 
    assign out[2790] = 1'b0; 
    assign out[2791] = 1'b0; 
    assign out[2792] = 1'b0; 
    assign out[2793] = 1'b0; 
    assign out[2794] = 1'b0; 
    assign out[2795] = 1'b0; 
    assign out[2796] = 1'b0; 
    assign out[2797] = 1'b0; 
    assign out[2798] = 1'b0; 
    assign out[2799] = 1'b0; 
    assign out[2800] = 1'b0; 
    assign out[2801] = 1'b0; 
    assign out[2802] = 1'b0; 
    assign out[2803] = 1'b0; 
    assign out[2804] = 1'b0; 
    assign out[2805] = 1'b0; 
    assign out[2806] = 1'b0; 
    assign out[2807] = 1'b0; 
    assign out[2808] = 1'b0; 
    assign out[2809] = 1'b0; 
    assign out[2810] = 1'b0; 
    assign out[2811] = 1'b0; 
    assign out[2812] = 1'b0; 
    assign out[2813] = 1'b0; 
    assign out[2814] = 1'b0; 
    assign out[2815] = 1'b0; 
    assign out[2816] = 1'b0; 
    assign out[2817] = 1'b0; 
    assign out[2818] = 1'b0; 
    assign out[2819] = 1'b0; 
    assign out[2820] = 1'b0; 
    assign out[2821] = 1'b0; 
    assign out[2822] = 1'b0; 
    assign out[2823] = 1'b0; 
    assign out[2824] = 1'b0; 
    assign out[2825] = 1'b0; 
    assign out[2826] = 1'b0; 
    assign out[2827] = 1'b0; 
    assign out[2828] = 1'b0; 
    assign out[2829] = 1'b0; 
    assign out[2830] = 1'b0; 
    assign out[2831] = 1'b0; 
    assign out[2832] = 1'b0; 
    assign out[2833] = 1'b0; 
    assign out[2834] = 1'b0; 
    assign out[2835] = 1'b0; 
    assign out[2836] = 1'b0; 
    assign out[2837] = 1'b0; 
    assign out[2838] = 1'b0; 
    assign out[2839] = 1'b0; 
    assign out[2840] = 1'b0; 
    assign out[2841] = 1'b0; 
    assign out[2842] = 1'b0; 
    assign out[2843] = 1'b0; 
    assign out[2844] = 1'b0; 
    assign out[2845] = 1'b0; 
    assign out[2846] = 1'b0; 
    assign out[2847] = 1'b0; 
    assign out[2848] = 1'b0; 
    assign out[2849] = 1'b0; 
    assign out[2850] = 1'b0; 
    assign out[2851] = 1'b0; 
    assign out[2852] = 1'b0; 
    assign out[2853] = 1'b0; 
    assign out[2854] = 1'b0; 
    assign out[2855] = 1'b0; 
    assign out[2856] = 1'b0; 
    assign out[2857] = 1'b0; 
    assign out[2858] = 1'b0; 
    assign out[2859] = 1'b0; 
    assign out[2860] = 1'b0; 
    assign out[2861] = 1'b0; 
    assign out[2862] = 1'b0; 
    assign out[2863] = 1'b0; 
    assign out[2864] = 1'b0; 
    assign out[2865] = 1'b0; 
    assign out[2866] = 1'b0; 
    assign out[2867] = 1'b0; 
    assign out[2868] = 1'b0; 
    assign out[2869] = 1'b0; 
    assign out[2870] = 1'b0; 
    assign out[2871] = 1'b0; 
    assign out[2872] = 1'b0; 
    assign out[2873] = 1'b0; 
    assign out[2874] = 1'b0; 
    assign out[2875] = 1'b0; 
    assign out[2876] = 1'b0; 
    assign out[2877] = 1'b0; 
    assign out[2878] = 1'b0; 
    assign out[2879] = 1'b0; 
    assign out[2880] = 1'b0; 
    assign out[2881] = 1'b0; 
    assign out[2882] = 1'b0; 
    assign out[2883] = 1'b0; 
    assign out[2884] = 1'b0; 
    assign out[2885] = 1'b0; 
    assign out[2886] = 1'b0; 
    assign out[2887] = 1'b0; 
    assign out[2888] = 1'b0; 
    assign out[2889] = 1'b0; 
    assign out[2890] = 1'b0; 
    assign out[2891] = 1'b0; 
    assign out[2892] = 1'b0; 
    assign out[2893] = 1'b0; 
    assign out[2894] = 1'b0; 
    assign out[2895] = 1'b0; 
    assign out[2896] = 1'b0; 
    assign out[2897] = 1'b0; 
    assign out[2898] = 1'b0; 
    assign out[2899] = 1'b0; 
    assign out[2900] = 1'b0; 
    assign out[2901] = 1'b0; 
    assign out[2902] = 1'b0; 
    assign out[2903] = 1'b0; 
    assign out[2904] = 1'b0; 
    assign out[2905] = 1'b0; 
    assign out[2906] = 1'b0; 
    assign out[2907] = 1'b0; 
    assign out[2908] = 1'b0; 
    assign out[2909] = 1'b0; 
    assign out[2910] = 1'b0; 
    assign out[2911] = 1'b0; 
    assign out[2912] = 1'b0; 
    assign out[2913] = 1'b0; 
    assign out[2914] = 1'b0; 
    assign out[2915] = 1'b0; 
    assign out[2916] = 1'b0; 
    assign out[2917] = 1'b0; 
    assign out[2918] = 1'b0; 
    assign out[2919] = 1'b0; 
    assign out[2920] = 1'b0; 
    assign out[2921] = 1'b0; 
    assign out[2922] = 1'b0; 
    assign out[2923] = 1'b0; 
    assign out[2924] = 1'b0; 
    assign out[2925] = 1'b0; 
    assign out[2926] = 1'b0; 
    assign out[2927] = 1'b0; 
    assign out[2928] = 1'b0; 
    assign out[2929] = 1'b0; 
    assign out[2930] = 1'b0; 
    assign out[2931] = 1'b0; 
    assign out[2932] = 1'b0; 
    assign out[2933] = 1'b0; 
    assign out[2934] = 1'b0; 
    assign out[2935] = 1'b0; 
    assign out[2936] = 1'b0; 
    assign out[2937] = 1'b0; 
    assign out[2938] = 1'b0; 
    assign out[2939] = 1'b0; 
    assign out[2940] = 1'b0; 
    assign out[2941] = 1'b0; 
    assign out[2942] = 1'b0; 
    assign out[2943] = 1'b0; 
    assign out[2944] = 1'b0; 
    assign out[2945] = 1'b0; 
    assign out[2946] = 1'b0; 
    assign out[2947] = 1'b0; 
    assign out[2948] = 1'b0; 
    assign out[2949] = 1'b0; 
    assign out[2950] = 1'b0; 
    assign out[2951] = 1'b0; 
    assign out[2952] = 1'b0; 
    assign out[2953] = 1'b0; 
    assign out[2954] = 1'b0; 
    assign out[2955] = 1'b0; 
    assign out[2956] = 1'b0; 
    assign out[2957] = 1'b0; 
    assign out[2958] = 1'b0; 
    assign out[2959] = 1'b0; 
    assign out[2960] = 1'b0; 
    assign out[2961] = 1'b0; 
    assign out[2962] = 1'b0; 
    assign out[2963] = 1'b0; 
    assign out[2964] = 1'b0; 
    assign out[2965] = 1'b0; 
    assign out[2966] = 1'b0; 
    assign out[2967] = 1'b0; 
    assign out[2968] = 1'b0; 
    assign out[2969] = 1'b0; 
    assign out[2970] = 1'b0; 
    assign out[2971] = 1'b0; 
    assign out[2972] = 1'b0; 
    assign out[2973] = 1'b0; 
    assign out[2974] = 1'b0; 
    assign out[2975] = 1'b0; 
    assign out[2976] = 1'b0; 
    assign out[2977] = 1'b0; 
    assign out[2978] = 1'b0; 
    assign out[2979] = 1'b0; 
    assign out[2980] = 1'b0; 
    assign out[2981] = 1'b0; 
    assign out[2982] = 1'b0; 
    assign out[2983] = 1'b0; 
    assign out[2984] = 1'b0; 
    assign out[2985] = 1'b0; 
    assign out[2986] = 1'b0; 
    assign out[2987] = 1'b0; 
    assign out[2988] = 1'b0; 
    assign out[2989] = 1'b0; 
    assign out[2990] = 1'b0; 
    assign out[2991] = 1'b0; 
    assign out[2992] = 1'b0; 
    assign out[2993] = 1'b0; 
    assign out[2994] = 1'b0; 
    assign out[2995] = 1'b0; 
    assign out[2996] = 1'b0; 
    assign out[2997] = 1'b0; 
    assign out[2998] = 1'b0; 
    assign out[2999] = 1'b0; 
    assign out[3000] = 1'b0; 
    assign out[3001] = 1'b0; 
    assign out[3002] = 1'b0; 
    assign out[3003] = 1'b0; 
    assign out[3004] = 1'b0; 
    assign out[3005] = 1'b0; 
    assign out[3006] = 1'b0; 
    assign out[3007] = 1'b0; 
    assign out[3008] = 1'b0; 
    assign out[3009] = 1'b0; 
    assign out[3010] = 1'b0; 
    assign out[3011] = 1'b0; 
    assign out[3012] = 1'b0; 
    assign out[3013] = 1'b0; 
    assign out[3014] = 1'b0; 
    assign out[3015] = 1'b0; 
    assign out[3016] = 1'b0; 
    assign out[3017] = 1'b0; 
    assign out[3018] = 1'b0; 
    assign out[3019] = 1'b0; 
    assign out[3020] = 1'b0; 
    assign out[3021] = 1'b0; 
    assign out[3022] = 1'b0; 
    assign out[3023] = 1'b0; 
    assign out[3024] = 1'b0; 
    assign out[3025] = 1'b0; 
    assign out[3026] = 1'b0; 
    assign out[3027] = 1'b0; 
    assign out[3028] = 1'b0; 
    assign out[3029] = 1'b0; 
    assign out[3030] = 1'b0; 
    assign out[3031] = 1'b0; 
    assign out[3032] = 1'b0; 
    assign out[3033] = 1'b0; 
    assign out[3034] = 1'b0; 
    assign out[3035] = 1'b0; 
    assign out[3036] = 1'b0; 
    assign out[3037] = 1'b0; 
    assign out[3038] = 1'b0; 
    assign out[3039] = 1'b0; 
    assign out[3040] = 1'b0; 
    assign out[3041] = 1'b0; 
    assign out[3042] = 1'b0; 
    assign out[3043] = 1'b0; 
    assign out[3044] = 1'b0; 
    assign out[3045] = 1'b0; 
    assign out[3046] = 1'b0; 
    assign out[3047] = 1'b0; 
    assign out[3048] = 1'b0; 
    assign out[3049] = 1'b0; 
    assign out[3050] = 1'b0; 
    assign out[3051] = 1'b0; 
    assign out[3052] = 1'b0; 
    assign out[3053] = 1'b0; 
    assign out[3054] = 1'b0; 
    assign out[3055] = 1'b0; 
    assign out[3056] = 1'b0; 
    assign out[3057] = 1'b0; 
    assign out[3058] = 1'b0; 
    assign out[3059] = 1'b0; 
    assign out[3060] = 1'b0; 
    assign out[3061] = 1'b0; 
    assign out[3062] = 1'b0; 
    assign out[3063] = 1'b0; 
    assign out[3064] = 1'b0; 
    assign out[3065] = 1'b0; 
    assign out[3066] = 1'b0; 
    assign out[3067] = 1'b0; 
    assign out[3068] = 1'b0; 
    assign out[3069] = 1'b0; 
    assign out[3070] = 1'b0; 
    assign out[3071] = 1'b0; 
    assign out[3072] = 1'b0; 
    assign out[3073] = 1'b0; 
    assign out[3074] = 1'b0; 
    assign out[3075] = 1'b0; 
    assign out[3076] = 1'b0; 
    assign out[3077] = 1'b0; 
    assign out[3078] = 1'b0; 
    assign out[3079] = 1'b0; 
    assign out[3080] = 1'b0; 
    assign out[3081] = 1'b0; 
    assign out[3082] = 1'b0; 
    assign out[3083] = 1'b0; 
    assign out[3084] = 1'b0; 
    assign out[3085] = 1'b0; 
    assign out[3086] = 1'b0; 
    assign out[3087] = 1'b0; 
    assign out[3088] = 1'b0; 
    assign out[3089] = 1'b0; 
    assign out[3090] = 1'b0; 
    assign out[3091] = 1'b0; 
    assign out[3092] = 1'b0; 
    assign out[3093] = 1'b0; 
    assign out[3094] = 1'b0; 
    assign out[3095] = 1'b0; 
    assign out[3096] = 1'b0; 
    assign out[3097] = 1'b0; 
    assign out[3098] = 1'b0; 
    assign out[3099] = 1'b0; 
    assign out[3100] = 1'b0; 
    assign out[3101] = 1'b0; 
    assign out[3102] = 1'b0; 
    assign out[3103] = 1'b0; 
    assign out[3104] = 1'b0; 
    assign out[3105] = 1'b0; 
    assign out[3106] = 1'b0; 
    assign out[3107] = 1'b0; 
    assign out[3108] = 1'b0; 
    assign out[3109] = 1'b0; 
    assign out[3110] = 1'b0; 
    assign out[3111] = 1'b0; 
    assign out[3112] = 1'b0; 
    assign out[3113] = 1'b0; 
    assign out[3114] = 1'b0; 
    assign out[3115] = 1'b0; 
    assign out[3116] = 1'b0; 
    assign out[3117] = 1'b0; 
    assign out[3118] = 1'b0; 
    assign out[3119] = 1'b0; 
    assign out[3120] = 1'b0; 
    assign out[3121] = 1'b0; 
    assign out[3122] = 1'b0; 
    assign out[3123] = 1'b0; 
    assign out[3124] = 1'b0; 
    assign out[3125] = 1'b0; 
    assign out[3126] = 1'b0; 
    assign out[3127] = 1'b0; 
    assign out[3128] = 1'b0; 
    assign out[3129] = 1'b0; 
    assign out[3130] = 1'b0; 
    assign out[3131] = 1'b0; 
    assign out[3132] = 1'b0; 
    assign out[3133] = 1'b0; 
    assign out[3134] = 1'b0; 
    assign out[3135] = 1'b0; 
    assign out[3136] = 1'b0; 
    assign out[3137] = 1'b0; 
    assign out[3138] = 1'b0; 
    assign out[3139] = 1'b0; 
    assign out[3140] = 1'b0; 
    assign out[3141] = 1'b0; 
    assign out[3142] = 1'b0; 
    assign out[3143] = 1'b0; 
    assign out[3144] = 1'b0; 
    assign out[3145] = 1'b0; 
    assign out[3146] = 1'b0; 
    assign out[3147] = 1'b0; 
    assign out[3148] = 1'b0; 
    assign out[3149] = 1'b0; 
    assign out[3150] = 1'b0; 
    assign out[3151] = 1'b0; 
    assign out[3152] = 1'b0; 
    assign out[3153] = 1'b0; 
    assign out[3154] = 1'b0; 
    assign out[3155] = 1'b0; 
    assign out[3156] = 1'b0; 
    assign out[3157] = 1'b0; 
    assign out[3158] = 1'b0; 
    assign out[3159] = 1'b0; 
    assign out[3160] = 1'b0; 
    assign out[3161] = 1'b0; 
    assign out[3162] = 1'b0; 
    assign out[3163] = 1'b0; 
    assign out[3164] = 1'b0; 
    assign out[3165] = 1'b0; 
    assign out[3166] = 1'b0; 
    assign out[3167] = 1'b0; 
    assign out[3168] = 1'b0; 
    assign out[3169] = 1'b0; 
    assign out[3170] = 1'b0; 
    assign out[3171] = 1'b0; 
    assign out[3172] = 1'b0; 
    assign out[3173] = 1'b0; 
    assign out[3174] = 1'b0; 
    assign out[3175] = 1'b0; 
    assign out[3176] = 1'b0; 
    assign out[3177] = 1'b0; 
    assign out[3178] = 1'b0; 
    assign out[3179] = 1'b0; 
    assign out[3180] = 1'b0; 
    assign out[3181] = 1'b0; 
    assign out[3182] = 1'b0; 
    assign out[3183] = 1'b0; 
    assign out[3184] = 1'b0; 
    assign out[3185] = 1'b0; 
    assign out[3186] = 1'b0; 
    assign out[3187] = 1'b0; 
    assign out[3188] = 1'b0; 
    assign out[3189] = 1'b0; 
    assign out[3190] = 1'b0; 
    assign out[3191] = 1'b0; 
    assign out[3192] = 1'b0; 
    assign out[3193] = 1'b0; 
    assign out[3194] = 1'b0; 
    assign out[3195] = 1'b0; 
    assign out[3196] = 1'b0; 
    assign out[3197] = 1'b0; 
    assign out[3198] = 1'b0; 
    assign out[3199] = 1'b0; 
    assign out[3200] = 1'b0; 
    assign out[3201] = 1'b0; 
    assign out[3202] = 1'b0; 
    assign out[3203] = 1'b0; 
    assign out[3204] = 1'b0; 
    assign out[3205] = 1'b0; 
    assign out[3206] = 1'b0; 
    assign out[3207] = 1'b0; 
    assign out[3208] = 1'b0; 
    assign out[3209] = 1'b0; 
    assign out[3210] = 1'b0; 
    assign out[3211] = 1'b0; 
    assign out[3212] = 1'b0; 
    assign out[3213] = 1'b0; 
    assign out[3214] = 1'b0; 
    assign out[3215] = 1'b0; 
    assign out[3216] = 1'b0; 
    assign out[3217] = 1'b0; 
    assign out[3218] = 1'b0; 
    assign out[3219] = 1'b0; 
    assign out[3220] = 1'b0; 
    assign out[3221] = 1'b0; 
    assign out[3222] = 1'b0; 
    assign out[3223] = 1'b0; 
    assign out[3224] = 1'b0; 
    assign out[3225] = 1'b0; 
    assign out[3226] = 1'b0; 
    assign out[3227] = 1'b0; 
    assign out[3228] = 1'b0; 
    assign out[3229] = 1'b0; 
    assign out[3230] = 1'b0; 
    assign out[3231] = 1'b0; 
    assign out[3232] = 1'b0; 
    assign out[3233] = 1'b0; 
    assign out[3234] = 1'b0; 
    assign out[3235] = 1'b0; 
    assign out[3236] = 1'b0; 
    assign out[3237] = 1'b0; 
    assign out[3238] = 1'b0; 
    assign out[3239] = 1'b0; 
    assign out[3240] = 1'b0; 
    assign out[3241] = 1'b0; 
    assign out[3242] = 1'b0; 
    assign out[3243] = 1'b0; 
    assign out[3244] = 1'b0; 
    assign out[3245] = 1'b0; 
    assign out[3246] = 1'b0; 
    assign out[3247] = 1'b0; 
    assign out[3248] = 1'b0; 
    assign out[3249] = 1'b0; 
    assign out[3250] = 1'b0; 
    assign out[3251] = 1'b0; 
    assign out[3252] = 1'b0; 
    assign out[3253] = 1'b0; 
    assign out[3254] = 1'b0; 
    assign out[3255] = 1'b0; 
    assign out[3256] = 1'b0; 
    assign out[3257] = 1'b0; 
    assign out[3258] = 1'b0; 
    assign out[3259] = 1'b0; 
    assign out[3260] = 1'b0; 
    assign out[3261] = 1'b0; 
    assign out[3262] = 1'b0; 
    assign out[3263] = 1'b0; 
    assign out[3264] = 1'b0; 
    assign out[3265] = 1'b0; 
    assign out[3266] = 1'b0; 
    assign out[3267] = 1'b0; 
    assign out[3268] = 1'b0; 
    assign out[3269] = 1'b0; 
    assign out[3270] = 1'b0; 
    assign out[3271] = 1'b0; 
    assign out[3272] = 1'b0; 
    assign out[3273] = 1'b0; 
    assign out[3274] = 1'b0; 
    assign out[3275] = 1'b0; 
    assign out[3276] = 1'b0; 
    assign out[3277] = 1'b0; 
    assign out[3278] = 1'b0; 
    assign out[3279] = 1'b0; 
    assign out[3280] = 1'b0; 
    assign out[3281] = 1'b0; 
    assign out[3282] = 1'b0; 
    assign out[3283] = 1'b0; 
    assign out[3284] = 1'b0; 
    assign out[3285] = 1'b0; 
    assign out[3286] = 1'b0; 
    assign out[3287] = 1'b0; 
    assign out[3288] = 1'b0; 
    assign out[3289] = 1'b0; 
    assign out[3290] = 1'b0; 
    assign out[3291] = 1'b0; 
    assign out[3292] = 1'b0; 
    assign out[3293] = 1'b0; 
    assign out[3294] = 1'b0; 
    assign out[3295] = 1'b0; 
    assign out[3296] = 1'b0; 
    assign out[3297] = 1'b0; 
    assign out[3298] = 1'b0; 
    assign out[3299] = 1'b0; 
    assign out[3300] = 1'b0; 
    assign out[3301] = 1'b0; 
    assign out[3302] = 1'b0; 
    assign out[3303] = 1'b0; 
    assign out[3304] = 1'b0; 
    assign out[3305] = 1'b0; 
    assign out[3306] = 1'b0; 
    assign out[3307] = 1'b0; 
    assign out[3308] = 1'b0; 
    assign out[3309] = 1'b0; 
    assign out[3310] = 1'b0; 
    assign out[3311] = 1'b0; 
    assign out[3312] = 1'b0; 
    assign out[3313] = 1'b0; 
    assign out[3314] = 1'b0; 
    assign out[3315] = 1'b0; 
    assign out[3316] = 1'b0; 
    assign out[3317] = 1'b0; 
    assign out[3318] = 1'b0; 
    assign out[3319] = 1'b0; 
    assign out[3320] = 1'b0; 
    assign out[3321] = 1'b0; 
    assign out[3322] = 1'b0; 
    assign out[3323] = 1'b0; 
    assign out[3324] = 1'b0; 
    assign out[3325] = 1'b0; 
    assign out[3326] = 1'b0; 
    assign out[3327] = 1'b0; 
    assign out[3328] = 1'b0; 
    assign out[3329] = 1'b0; 
    assign out[3330] = 1'b0; 
    assign out[3331] = 1'b0; 
    assign out[3332] = 1'b0; 
    assign out[3333] = 1'b0; 
    assign out[3334] = 1'b0; 
    assign out[3335] = 1'b0; 
    assign out[3336] = 1'b0; 
    assign out[3337] = 1'b0; 
    assign out[3338] = 1'b0; 
    assign out[3339] = 1'b0; 
    assign out[3340] = 1'b0; 
    assign out[3341] = 1'b0; 
    assign out[3342] = 1'b0; 
    assign out[3343] = 1'b0; 
    assign out[3344] = 1'b0; 
    assign out[3345] = 1'b0; 
    assign out[3346] = 1'b0; 
    assign out[3347] = 1'b0; 
    assign out[3348] = 1'b0; 
    assign out[3349] = 1'b0; 
    assign out[3350] = 1'b0; 
    assign out[3351] = 1'b0; 
    assign out[3352] = 1'b0; 
    assign out[3353] = 1'b0; 
    assign out[3354] = 1'b0; 
    assign out[3355] = 1'b0; 
    assign out[3356] = 1'b0; 
    assign out[3357] = 1'b0; 
    assign out[3358] = 1'b0; 
    assign out[3359] = 1'b0; 
    assign out[3360] = 1'b0; 
    assign out[3361] = 1'b0; 
    assign out[3362] = 1'b0; 
    assign out[3363] = 1'b0; 
    assign out[3364] = 1'b0; 
    assign out[3365] = 1'b0; 
    assign out[3366] = 1'b0; 
    assign out[3367] = 1'b0; 
    assign out[3368] = 1'b0; 
    assign out[3369] = 1'b0; 
    assign out[3370] = 1'b0; 
    assign out[3371] = 1'b0; 
    assign out[3372] = 1'b0; 
    assign out[3373] = 1'b0; 
    assign out[3374] = 1'b0; 
    assign out[3375] = 1'b0; 
    assign out[3376] = 1'b0; 
    assign out[3377] = 1'b0; 
    assign out[3378] = 1'b0; 
    assign out[3379] = 1'b0; 
    assign out[3380] = 1'b0; 
    assign out[3381] = 1'b0; 
    assign out[3382] = 1'b0; 
    assign out[3383] = 1'b0; 
    assign out[3384] = 1'b0; 
    assign out[3385] = 1'b0; 
    assign out[3386] = 1'b0; 
    assign out[3387] = 1'b0; 
    assign out[3388] = 1'b0; 
    assign out[3389] = 1'b0; 
    assign out[3390] = 1'b0; 
    assign out[3391] = 1'b0; 
    assign out[3392] = 1'b0; 
    assign out[3393] = 1'b0; 
    assign out[3394] = 1'b0; 
    assign out[3395] = 1'b0; 
    assign out[3396] = 1'b0; 
    assign out[3397] = 1'b0; 
    assign out[3398] = 1'b0; 
    assign out[3399] = 1'b0; 
    assign out[3400] = 1'b0; 
    assign out[3401] = 1'b0; 
    assign out[3402] = 1'b0; 
    assign out[3403] = 1'b0; 
    assign out[3404] = 1'b0; 
    assign out[3405] = 1'b0; 
    assign out[3406] = 1'b0; 
    assign out[3407] = 1'b0; 
    assign out[3408] = 1'b0; 
    assign out[3409] = 1'b0; 
    assign out[3410] = 1'b0; 
    assign out[3411] = 1'b0; 
    assign out[3412] = 1'b0; 
    assign out[3413] = 1'b0; 
    assign out[3414] = 1'b0; 
    assign out[3415] = 1'b0; 
    assign out[3416] = 1'b0; 
    assign out[3417] = 1'b0; 
    assign out[3418] = 1'b0; 
    assign out[3419] = 1'b0; 
    assign out[3420] = 1'b0; 
    assign out[3421] = 1'b0; 
    assign out[3422] = 1'b0; 
    assign out[3423] = 1'b0; 
    assign out[3424] = 1'b0; 
    assign out[3425] = 1'b0; 
    assign out[3426] = 1'b0; 
    assign out[3427] = 1'b0; 
    assign out[3428] = 1'b0; 
    assign out[3429] = 1'b0; 
    assign out[3430] = 1'b0; 
    assign out[3431] = 1'b0; 
    assign out[3432] = 1'b0; 
    assign out[3433] = 1'b0; 
    assign out[3434] = 1'b0; 
    assign out[3435] = 1'b0; 
    assign out[3436] = 1'b0; 
    assign out[3437] = 1'b0; 
    assign out[3438] = 1'b0; 
    assign out[3439] = 1'b0; 
    assign out[3440] = 1'b0; 
    assign out[3441] = 1'b0; 
    assign out[3442] = 1'b0; 
    assign out[3443] = 1'b0; 
    assign out[3444] = 1'b0; 
    assign out[3445] = 1'b0; 
    assign out[3446] = 1'b0; 
    assign out[3447] = 1'b0; 
    assign out[3448] = 1'b0; 
    assign out[3449] = 1'b0; 
    assign out[3450] = 1'b0; 
    assign out[3451] = 1'b0; 
    assign out[3452] = 1'b0; 
    assign out[3453] = 1'b0; 
    assign out[3454] = 1'b0; 
    assign out[3455] = 1'b0; 
    assign out[3456] = 1'b0; 
    assign out[3457] = 1'b0; 
    assign out[3458] = 1'b0; 
    assign out[3459] = 1'b0; 
    assign out[3460] = 1'b0; 
    assign out[3461] = 1'b0; 
    assign out[3462] = 1'b0; 
    assign out[3463] = 1'b0; 
    assign out[3464] = 1'b0; 
    assign out[3465] = 1'b0; 
    assign out[3466] = 1'b0; 
    assign out[3467] = 1'b0; 
    assign out[3468] = 1'b0; 
    assign out[3469] = 1'b0; 
    assign out[3470] = 1'b0; 
    assign out[3471] = 1'b0; 
    assign out[3472] = 1'b0; 
    assign out[3473] = 1'b0; 
    assign out[3474] = 1'b0; 
    assign out[3475] = 1'b0; 
    assign out[3476] = 1'b0; 
    assign out[3477] = 1'b0; 
    assign out[3478] = 1'b0; 
    assign out[3479] = 1'b0; 
    assign out[3480] = 1'b0; 
    assign out[3481] = 1'b0; 
    assign out[3482] = 1'b0; 
    assign out[3483] = 1'b0; 
    assign out[3484] = 1'b0; 
    assign out[3485] = 1'b0; 
    assign out[3486] = 1'b0; 
    assign out[3487] = 1'b0; 
    assign out[3488] = 1'b0; 
    assign out[3489] = 1'b0; 
    assign out[3490] = 1'b0; 
    assign out[3491] = 1'b0; 
    assign out[3492] = 1'b0; 
    assign out[3493] = 1'b0; 
    assign out[3494] = 1'b0; 
    assign out[3495] = 1'b0; 
    assign out[3496] = 1'b0; 
    assign out[3497] = 1'b0; 
    assign out[3498] = 1'b0; 
    assign out[3499] = 1'b0; 
    assign out[3500] = 1'b0; 
    assign out[3501] = 1'b0; 
    assign out[3502] = 1'b0; 
    assign out[3503] = 1'b0; 
    assign out[3504] = 1'b0; 
    assign out[3505] = 1'b0; 
    assign out[3506] = 1'b0; 
    assign out[3507] = 1'b0; 
    assign out[3508] = 1'b0; 
    assign out[3509] = 1'b0; 
    assign out[3510] = 1'b0; 
    assign out[3511] = 1'b0; 
    assign out[3512] = 1'b0; 
    assign out[3513] = 1'b0; 
    assign out[3514] = 1'b0; 
    assign out[3515] = 1'b0; 
    assign out[3516] = 1'b0; 
    assign out[3517] = 1'b0; 
    assign out[3518] = 1'b0; 
    assign out[3519] = 1'b0; 
    assign out[3520] = 1'b0; 
    assign out[3521] = 1'b0; 
    assign out[3522] = 1'b0; 
    assign out[3523] = 1'b0; 
    assign out[3524] = 1'b0; 
    assign out[3525] = 1'b0; 
    assign out[3526] = 1'b0; 
    assign out[3527] = 1'b0; 
    assign out[3528] = 1'b0; 
    assign out[3529] = 1'b0; 
    assign out[3530] = 1'b0; 
    assign out[3531] = 1'b0; 
    assign out[3532] = 1'b0; 
    assign out[3533] = 1'b0; 
    assign out[3534] = 1'b0; 
    assign out[3535] = 1'b0; 
    assign out[3536] = 1'b0; 
    assign out[3537] = 1'b0; 
    assign out[3538] = 1'b0; 
    assign out[3539] = 1'b0; 
    assign out[3540] = 1'b0; 
    assign out[3541] = 1'b0; 
    assign out[3542] = 1'b0; 
    assign out[3543] = 1'b0; 
    assign out[3544] = 1'b0; 
    assign out[3545] = 1'b0; 
    assign out[3546] = 1'b0; 
    assign out[3547] = 1'b0; 
    assign out[3548] = 1'b0; 
    assign out[3549] = 1'b0; 
    assign out[3550] = 1'b0; 
    assign out[3551] = 1'b0; 
    assign out[3552] = 1'b0; 
    assign out[3553] = 1'b0; 
    assign out[3554] = 1'b0; 
    assign out[3555] = 1'b0; 
    assign out[3556] = 1'b0; 
    assign out[3557] = 1'b0; 
    assign out[3558] = 1'b0; 
    assign out[3559] = 1'b0; 
    assign out[3560] = 1'b0; 
    assign out[3561] = 1'b0; 
    assign out[3562] = 1'b0; 
    assign out[3563] = 1'b0; 
    assign out[3564] = 1'b0; 
    assign out[3565] = 1'b0; 
    assign out[3566] = 1'b0; 
    assign out[3567] = 1'b0; 
    assign out[3568] = 1'b0; 
    assign out[3569] = 1'b0; 
    assign out[3570] = 1'b0; 
    assign out[3571] = 1'b0; 
    assign out[3572] = 1'b0; 
    assign out[3573] = 1'b0; 
    assign out[3574] = 1'b0; 
    assign out[3575] = 1'b0; 
    assign out[3576] = 1'b0; 
    assign out[3577] = 1'b0; 
    assign out[3578] = 1'b0; 
    assign out[3579] = 1'b0; 
    assign out[3580] = 1'b0; 
    assign out[3581] = 1'b0; 
    assign out[3582] = 1'b0; 
    assign out[3583] = 1'b0; 
    assign out[3584] = 1'b0; 
    assign out[3585] = 1'b0; 
    assign out[3586] = 1'b0; 
    assign out[3587] = 1'b0; 
    assign out[3588] = 1'b0; 
    assign out[3589] = 1'b0; 
    assign out[3590] = 1'b0; 
    assign out[3591] = 1'b0; 
    assign out[3592] = 1'b0; 
    assign out[3593] = 1'b0; 
    assign out[3594] = 1'b0; 
    assign out[3595] = 1'b0; 
    assign out[3596] = 1'b0; 
    assign out[3597] = 1'b0; 
    assign out[3598] = 1'b0; 
    assign out[3599] = 1'b0; 
    assign out[3600] = 1'b0; 
    assign out[3601] = 1'b0; 
    assign out[3602] = 1'b0; 
    assign out[3603] = 1'b0; 
    assign out[3604] = 1'b0; 
    assign out[3605] = 1'b0; 
    assign out[3606] = 1'b0; 
    assign out[3607] = 1'b0; 
    assign out[3608] = 1'b0; 
    assign out[3609] = 1'b0; 
    assign out[3610] = 1'b0; 
    assign out[3611] = 1'b0; 
    assign out[3612] = 1'b0; 
    assign out[3613] = 1'b0; 
    assign out[3614] = 1'b0; 
    assign out[3615] = 1'b0; 
    assign out[3616] = 1'b0; 
    assign out[3617] = 1'b0; 
    assign out[3618] = 1'b0; 
    assign out[3619] = 1'b0; 
    assign out[3620] = 1'b0; 
    assign out[3621] = 1'b0; 
    assign out[3622] = 1'b0; 
    assign out[3623] = 1'b0; 
    assign out[3624] = 1'b0; 
    assign out[3625] = 1'b0; 
    assign out[3626] = 1'b0; 
    assign out[3627] = 1'b0; 
    assign out[3628] = 1'b0; 
    assign out[3629] = 1'b0; 
    assign out[3630] = 1'b0; 
    assign out[3631] = 1'b0; 
    assign out[3632] = 1'b0; 
    assign out[3633] = 1'b0; 
    assign out[3634] = 1'b0; 
    assign out[3635] = 1'b0; 
    assign out[3636] = 1'b0; 
    assign out[3637] = 1'b0; 
    assign out[3638] = 1'b0; 
    assign out[3639] = 1'b0; 
    assign out[3640] = 1'b0; 
    assign out[3641] = 1'b0; 
    assign out[3642] = 1'b0; 
    assign out[3643] = 1'b0; 
    assign out[3644] = 1'b0; 
    assign out[3645] = 1'b0; 
    assign out[3646] = 1'b0; 
    assign out[3647] = 1'b0; 
    assign out[3648] = 1'b0; 
    assign out[3649] = 1'b0; 
    assign out[3650] = 1'b0; 
    assign out[3651] = 1'b0; 
    assign out[3652] = 1'b0; 
    assign out[3653] = 1'b0; 
    assign out[3654] = 1'b0; 
    assign out[3655] = 1'b0; 
    assign out[3656] = 1'b0; 
    assign out[3657] = 1'b0; 
    assign out[3658] = 1'b0; 
    assign out[3659] = 1'b0; 
    assign out[3660] = 1'b0; 
    assign out[3661] = 1'b0; 
    assign out[3662] = 1'b0; 
    assign out[3663] = 1'b0; 
    assign out[3664] = 1'b0; 
    assign out[3665] = 1'b0; 
    assign out[3666] = 1'b0; 
    assign out[3667] = 1'b0; 
    assign out[3668] = 1'b0; 
    assign out[3669] = 1'b0; 
    assign out[3670] = 1'b0; 
    assign out[3671] = 1'b0; 
    assign out[3672] = 1'b0; 
    assign out[3673] = 1'b0; 
    assign out[3674] = 1'b0; 
    assign out[3675] = 1'b0; 
    assign out[3676] = 1'b0; 
    assign out[3677] = 1'b0; 
    assign out[3678] = 1'b0; 
    assign out[3679] = 1'b0; 
    assign out[3680] = 1'b0; 
    assign out[3681] = 1'b0; 
    assign out[3682] = 1'b0; 
    assign out[3683] = 1'b0; 
    assign out[3684] = 1'b0; 
    assign out[3685] = 1'b0; 
    assign out[3686] = 1'b0; 
    assign out[3687] = 1'b0; 
    assign out[3688] = 1'b0; 
    assign out[3689] = 1'b0; 
    assign out[3690] = 1'b0; 
    assign out[3691] = 1'b0; 
    assign out[3692] = 1'b0; 
    assign out[3693] = 1'b0; 
    assign out[3694] = 1'b0; 
    assign out[3695] = 1'b0; 
    assign out[3696] = 1'b0; 
    assign out[3697] = 1'b0; 
    assign out[3698] = 1'b0; 
    assign out[3699] = 1'b0; 
    assign out[3700] = 1'b0; 
    assign out[3701] = 1'b0; 
    assign out[3702] = 1'b0; 
    assign out[3703] = 1'b0; 
    assign out[3704] = 1'b0; 
    assign out[3705] = 1'b0; 
    assign out[3706] = 1'b0; 
    assign out[3707] = 1'b0; 
    assign out[3708] = 1'b0; 
    assign out[3709] = 1'b0; 
    assign out[3710] = 1'b0; 
    assign out[3711] = 1'b0; 
    assign out[3712] = 1'b0; 
    assign out[3713] = 1'b0; 
    assign out[3714] = 1'b0; 
    assign out[3715] = 1'b0; 
    assign out[3716] = 1'b0; 
    assign out[3717] = 1'b0; 
    assign out[3718] = 1'b0; 
    assign out[3719] = 1'b0; 
    assign out[3720] = 1'b0; 
    assign out[3721] = 1'b0; 
    assign out[3722] = 1'b0; 
    assign out[3723] = 1'b0; 
    assign out[3724] = 1'b0; 
    assign out[3725] = 1'b0; 
    assign out[3726] = 1'b0; 
    assign out[3727] = 1'b0; 
    assign out[3728] = 1'b0; 
    assign out[3729] = 1'b0; 
    assign out[3730] = 1'b0; 
    assign out[3731] = 1'b0; 
    assign out[3732] = 1'b0; 
    assign out[3733] = 1'b0; 
    assign out[3734] = 1'b0; 
    assign out[3735] = 1'b0; 
    assign out[3736] = 1'b0; 
    assign out[3737] = 1'b0; 
    assign out[3738] = 1'b0; 
    assign out[3739] = 1'b0; 
    assign out[3740] = 1'b0; 
    assign out[3741] = 1'b0; 
    assign out[3742] = 1'b0; 
    assign out[3743] = 1'b0; 
    assign out[3744] = 1'b0; 
    assign out[3745] = 1'b0; 
    assign out[3746] = 1'b0; 
    assign out[3747] = 1'b0; 
    assign out[3748] = 1'b0; 
    assign out[3749] = 1'b0; 
    assign out[3750] = 1'b0; 
    assign out[3751] = 1'b0; 
    assign out[3752] = 1'b0; 
    assign out[3753] = 1'b0; 
    assign out[3754] = 1'b0; 
    assign out[3755] = 1'b0; 
    assign out[3756] = 1'b0; 
    assign out[3757] = 1'b0; 
    assign out[3758] = 1'b0; 
    assign out[3759] = 1'b0; 
    assign out[3760] = 1'b0; 
    assign out[3761] = 1'b0; 
    assign out[3762] = 1'b0; 
    assign out[3763] = 1'b0; 
    assign out[3764] = 1'b0; 
    assign out[3765] = 1'b0; 
    assign out[3766] = 1'b0; 
    assign out[3767] = 1'b0; 
    assign out[3768] = 1'b0; 
    assign out[3769] = 1'b0; 
    assign out[3770] = 1'b0; 
    assign out[3771] = 1'b0; 
    assign out[3772] = 1'b0; 
    assign out[3773] = 1'b0; 
    assign out[3774] = 1'b0; 
    assign out[3775] = 1'b0; 
    assign out[3776] = 1'b0; 
    assign out[3777] = 1'b0; 
    assign out[3778] = 1'b0; 
    assign out[3779] = 1'b0; 
    assign out[3780] = 1'b0; 
    assign out[3781] = 1'b0; 
    assign out[3782] = 1'b0; 
    assign out[3783] = 1'b0; 
    assign out[3784] = 1'b0; 
    assign out[3785] = 1'b0; 
    assign out[3786] = 1'b0; 
    assign out[3787] = 1'b0; 
    assign out[3788] = 1'b0; 
    assign out[3789] = 1'b0; 
    assign out[3790] = 1'b0; 
    assign out[3791] = 1'b0; 
    assign out[3792] = 1'b0; 
    assign out[3793] = 1'b0; 
    assign out[3794] = 1'b0; 
    assign out[3795] = 1'b0; 
    assign out[3796] = 1'b0; 
    assign out[3797] = 1'b0; 
    assign out[3798] = 1'b0; 
    assign out[3799] = 1'b0; 
    assign out[3800] = 1'b0; 
    assign out[3801] = 1'b0; 
    assign out[3802] = 1'b0; 
    assign out[3803] = 1'b0; 
    assign out[3804] = 1'b0; 
    assign out[3805] = 1'b0; 
    assign out[3806] = 1'b0; 
    assign out[3807] = 1'b0; 
    assign out[3808] = 1'b0; 
    assign out[3809] = 1'b0; 
    assign out[3810] = 1'b0; 
    assign out[3811] = 1'b0; 
    assign out[3812] = 1'b0; 
    assign out[3813] = 1'b0; 
    assign out[3814] = 1'b0; 
    assign out[3815] = 1'b0; 
    assign out[3816] = 1'b0; 
    assign out[3817] = 1'b0; 
    assign out[3818] = 1'b0; 
    assign out[3819] = 1'b0; 
    assign out[3820] = 1'b0; 
    assign out[3821] = 1'b0; 
    assign out[3822] = 1'b0; 
    assign out[3823] = 1'b0; 
    assign out[3824] = 1'b0; 
    assign out[3825] = 1'b0; 
    assign out[3826] = 1'b0; 
    assign out[3827] = 1'b0; 
    assign out[3828] = 1'b0; 
    assign out[3829] = 1'b0; 
    assign out[3830] = 1'b0; 
    assign out[3831] = 1'b0; 
    assign out[3832] = 1'b0; 
    assign out[3833] = 1'b0; 
    assign out[3834] = 1'b0; 
    assign out[3835] = 1'b0; 
    assign out[3836] = 1'b0; 
    assign out[3837] = 1'b0; 
    assign out[3838] = 1'b0; 
    assign out[3839] = 1'b0; 
    assign out[3840] = 1'b0; 
    assign out[3841] = 1'b0; 
    assign out[3842] = 1'b0; 
    assign out[3843] = 1'b0; 
    assign out[3844] = 1'b0; 
    assign out[3845] = 1'b0; 
    assign out[3846] = 1'b0; 
    assign out[3847] = 1'b0; 
    assign out[3848] = 1'b0; 
    assign out[3849] = 1'b0; 
    assign out[3850] = 1'b0; 
    assign out[3851] = 1'b0; 
    assign out[3852] = 1'b0; 
    assign out[3853] = 1'b0; 
    assign out[3854] = 1'b0; 
    assign out[3855] = 1'b0; 
    assign out[3856] = 1'b0; 
    assign out[3857] = 1'b0; 
    assign out[3858] = 1'b0; 
    assign out[3859] = 1'b0; 
    assign out[3860] = 1'b0; 
    assign out[3861] = 1'b0; 
    assign out[3862] = 1'b0; 
    assign out[3863] = 1'b0; 
    assign out[3864] = 1'b0; 
    assign out[3865] = 1'b0; 
    assign out[3866] = 1'b0; 
    assign out[3867] = 1'b0; 
    assign out[3868] = 1'b0; 
    assign out[3869] = 1'b0; 
    assign out[3870] = 1'b0; 
    assign out[3871] = 1'b0; 
    assign out[3872] = 1'b0; 
    assign out[3873] = 1'b0; 
    assign out[3874] = 1'b0; 
    assign out[3875] = 1'b0; 
    assign out[3876] = 1'b0; 
    assign out[3877] = 1'b0; 
    assign out[3878] = 1'b0; 
    assign out[3879] = 1'b0; 
    assign out[3880] = 1'b0; 
    assign out[3881] = 1'b0; 
    assign out[3882] = 1'b0; 
    assign out[3883] = 1'b0; 
    assign out[3884] = 1'b0; 
    assign out[3885] = 1'b0; 
    assign out[3886] = 1'b0; 
    assign out[3887] = 1'b0; 
    assign out[3888] = 1'b0; 
    assign out[3889] = 1'b0; 
    assign out[3890] = 1'b0; 
    assign out[3891] = 1'b0; 
    assign out[3892] = 1'b0; 
    assign out[3893] = 1'b0; 
    assign out[3894] = 1'b0; 
    assign out[3895] = 1'b0; 
    assign out[3896] = 1'b0; 
    assign out[3897] = 1'b0; 
    assign out[3898] = 1'b0; 
    assign out[3899] = 1'b0; 
    assign out[3900] = 1'b0; 
    assign out[3901] = 1'b0; 
    assign out[3902] = 1'b0; 
    assign out[3903] = 1'b0; 
    assign out[3904] = 1'b0; 
    assign out[3905] = 1'b0; 
    assign out[3906] = 1'b0; 
    assign out[3907] = 1'b0; 
    assign out[3908] = 1'b0; 
    assign out[3909] = 1'b0; 
    assign out[3910] = 1'b0; 
    assign out[3911] = 1'b0; 
    assign out[3912] = 1'b0; 
    assign out[3913] = 1'b0; 
    assign out[3914] = 1'b0; 
    assign out[3915] = 1'b0; 
    assign out[3916] = 1'b0; 
    assign out[3917] = 1'b0; 
    assign out[3918] = 1'b0; 
    assign out[3919] = 1'b0; 
    assign out[3920] = 1'b0; 
    assign out[3921] = 1'b0; 
    assign out[3922] = 1'b0; 
    assign out[3923] = 1'b0; 
    assign out[3924] = 1'b0; 
    assign out[3925] = 1'b0; 
    assign out[3926] = 1'b0; 
    assign out[3927] = 1'b0; 
    assign out[3928] = 1'b0; 
    assign out[3929] = 1'b0; 
    assign out[3930] = 1'b0; 
    assign out[3931] = 1'b0; 
    assign out[3932] = 1'b0; 
    assign out[3933] = 1'b0; 
    assign out[3934] = 1'b0; 
    assign out[3935] = 1'b0; 
    assign out[3936] = 1'b0; 
    assign out[3937] = 1'b0; 
    assign out[3938] = 1'b0; 
    assign out[3939] = 1'b0; 
    assign out[3940] = 1'b0; 
    assign out[3941] = 1'b0; 
    assign out[3942] = 1'b0; 
    assign out[3943] = 1'b0; 
    assign out[3944] = 1'b0; 
    assign out[3945] = 1'b0; 
    assign out[3946] = 1'b0; 
    assign out[3947] = 1'b0; 
    assign out[3948] = 1'b0; 
    assign out[3949] = 1'b0; 
    assign out[3950] = 1'b0; 
    assign out[3951] = 1'b0; 
    assign out[3952] = 1'b0; 
    assign out[3953] = 1'b0; 
    assign out[3954] = 1'b0; 
    assign out[3955] = 1'b0; 
    assign out[3956] = 1'b0; 
    assign out[3957] = 1'b0; 
    assign out[3958] = 1'b0; 
    assign out[3959] = 1'b0; 
    assign out[3960] = 1'b0; 
    assign out[3961] = 1'b0; 
    assign out[3962] = 1'b0; 
    assign out[3963] = 1'b0; 
    assign out[3964] = 1'b0; 
    assign out[3965] = 1'b0; 
    assign out[3966] = 1'b0; 
    assign out[3967] = 1'b0; 
    assign out[3968] = 1'b0; 
    assign out[3969] = 1'b0; 
    assign out[3970] = 1'b0; 
    assign out[3971] = 1'b0; 
    assign out[3972] = 1'b0; 
    assign out[3973] = 1'b0; 
    assign out[3974] = 1'b0; 
    assign out[3975] = 1'b0; 
    assign out[3976] = 1'b0; 
    assign out[3977] = 1'b0; 
    assign out[3978] = 1'b0; 
    assign out[3979] = 1'b0; 
    assign out[3980] = 1'b0; 
    assign out[3981] = 1'b0; 
    assign out[3982] = 1'b0; 
    assign out[3983] = 1'b0; 
    assign out[3984] = 1'b0; 
    assign out[3985] = 1'b0; 
    assign out[3986] = 1'b0; 
    assign out[3987] = 1'b0; 
    assign out[3988] = 1'b0; 
    assign out[3989] = 1'b0; 
    assign out[3990] = 1'b0; 
    assign out[3991] = 1'b0; 
    assign out[3992] = 1'b0; 
    assign out[3993] = 1'b0; 
    assign out[3994] = 1'b0; 
    assign out[3995] = 1'b0; 
    assign out[3996] = 1'b0; 
    assign out[3997] = 1'b0; 
    assign out[3998] = 1'b0; 
    assign out[3999] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[2549:0] = out[2549:0];

endmodule
