magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -696 -419 696 419
<< pmos >>
rect -500 -200 500 200
<< pdiff >>
rect -558 187 -500 200
rect -558 153 -546 187
rect -512 153 -500 187
rect -558 119 -500 153
rect -558 85 -546 119
rect -512 85 -500 119
rect -558 51 -500 85
rect -558 17 -546 51
rect -512 17 -500 51
rect -558 -17 -500 17
rect -558 -51 -546 -17
rect -512 -51 -500 -17
rect -558 -85 -500 -51
rect -558 -119 -546 -85
rect -512 -119 -500 -85
rect -558 -153 -500 -119
rect -558 -187 -546 -153
rect -512 -187 -500 -153
rect -558 -200 -500 -187
rect 500 187 558 200
rect 500 153 512 187
rect 546 153 558 187
rect 500 119 558 153
rect 500 85 512 119
rect 546 85 558 119
rect 500 51 558 85
rect 500 17 512 51
rect 546 17 558 51
rect 500 -17 558 17
rect 500 -51 512 -17
rect 546 -51 558 -17
rect 500 -85 558 -51
rect 500 -119 512 -85
rect 546 -119 558 -85
rect 500 -153 558 -119
rect 500 -187 512 -153
rect 546 -187 558 -153
rect 500 -200 558 -187
<< pdiffc >>
rect -546 153 -512 187
rect -546 85 -512 119
rect -546 17 -512 51
rect -546 -51 -512 -17
rect -546 -119 -512 -85
rect -546 -187 -512 -153
rect 512 153 546 187
rect 512 85 546 119
rect 512 17 546 51
rect 512 -51 546 -17
rect 512 -119 546 -85
rect 512 -187 546 -153
<< nsubdiff >>
rect -660 349 -561 383
rect -527 349 -493 383
rect -459 349 -425 383
rect -391 349 -357 383
rect -323 349 -289 383
rect -255 349 -221 383
rect -187 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 187 383
rect 221 349 255 383
rect 289 349 323 383
rect 357 349 391 383
rect 425 349 459 383
rect 493 349 527 383
rect 561 349 660 383
rect -660 255 -626 349
rect -660 187 -626 221
rect 626 255 660 349
rect -660 119 -626 153
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect -660 -153 -626 -119
rect -660 -221 -626 -187
rect 626 187 660 221
rect 626 119 660 153
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect 626 -153 660 -119
rect -660 -349 -626 -255
rect 626 -221 660 -187
rect 626 -349 660 -255
rect -660 -383 -561 -349
rect -527 -383 -493 -349
rect -459 -383 -425 -349
rect -391 -383 -357 -349
rect -323 -383 -289 -349
rect -255 -383 -221 -349
rect -187 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 187 -349
rect 221 -383 255 -349
rect 289 -383 323 -349
rect 357 -383 391 -349
rect 425 -383 459 -349
rect 493 -383 527 -349
rect 561 -383 660 -349
<< nsubdiffcont >>
rect -561 349 -527 383
rect -493 349 -459 383
rect -425 349 -391 383
rect -357 349 -323 383
rect -289 349 -255 383
rect -221 349 -187 383
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect 187 349 221 383
rect 255 349 289 383
rect 323 349 357 383
rect 391 349 425 383
rect 459 349 493 383
rect 527 349 561 383
rect -660 221 -626 255
rect 626 221 660 255
rect -660 153 -626 187
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -660 -187 -626 -153
rect 626 153 660 187
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect 626 -187 660 -153
rect -660 -255 -626 -221
rect 626 -255 660 -221
rect -561 -383 -527 -349
rect -493 -383 -459 -349
rect -425 -383 -391 -349
rect -357 -383 -323 -349
rect -289 -383 -255 -349
rect -221 -383 -187 -349
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
rect 187 -383 221 -349
rect 255 -383 289 -349
rect 323 -383 357 -349
rect 391 -383 425 -349
rect 459 -383 493 -349
rect 527 -383 561 -349
<< poly >>
rect -500 281 500 297
rect -500 247 -459 281
rect -425 247 -391 281
rect -357 247 -323 281
rect -289 247 -255 281
rect -221 247 -187 281
rect -153 247 -119 281
rect -85 247 -51 281
rect -17 247 17 281
rect 51 247 85 281
rect 119 247 153 281
rect 187 247 221 281
rect 255 247 289 281
rect 323 247 357 281
rect 391 247 425 281
rect 459 247 500 281
rect -500 200 500 247
rect -500 -247 500 -200
rect -500 -281 -459 -247
rect -425 -281 -391 -247
rect -357 -281 -323 -247
rect -289 -281 -255 -247
rect -221 -281 -187 -247
rect -153 -281 -119 -247
rect -85 -281 -51 -247
rect -17 -281 17 -247
rect 51 -281 85 -247
rect 119 -281 153 -247
rect 187 -281 221 -247
rect 255 -281 289 -247
rect 323 -281 357 -247
rect 391 -281 425 -247
rect 459 -281 500 -247
rect -500 -297 500 -281
<< polycont >>
rect -459 247 -425 281
rect -391 247 -357 281
rect -323 247 -289 281
rect -255 247 -221 281
rect -187 247 -153 281
rect -119 247 -85 281
rect -51 247 -17 281
rect 17 247 51 281
rect 85 247 119 281
rect 153 247 187 281
rect 221 247 255 281
rect 289 247 323 281
rect 357 247 391 281
rect 425 247 459 281
rect -459 -281 -425 -247
rect -391 -281 -357 -247
rect -323 -281 -289 -247
rect -255 -281 -221 -247
rect -187 -281 -153 -247
rect -119 -281 -85 -247
rect -51 -281 -17 -247
rect 17 -281 51 -247
rect 85 -281 119 -247
rect 153 -281 187 -247
rect 221 -281 255 -247
rect 289 -281 323 -247
rect 357 -281 391 -247
rect 425 -281 459 -247
<< locali >>
rect -660 349 -561 383
rect -527 349 -493 383
rect -459 349 -425 383
rect -391 349 -357 383
rect -323 349 -289 383
rect -255 349 -221 383
rect -187 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 187 383
rect 221 349 255 383
rect 289 349 323 383
rect 357 349 391 383
rect 425 349 459 383
rect 493 349 527 383
rect 561 349 660 383
rect -660 255 -626 349
rect -500 247 -459 281
rect -415 247 -391 281
rect -343 247 -323 281
rect -271 247 -255 281
rect -199 247 -187 281
rect -127 247 -119 281
rect -55 247 -51 281
rect 51 247 55 281
rect 119 247 127 281
rect 187 247 199 281
rect 255 247 271 281
rect 323 247 343 281
rect 391 247 415 281
rect 459 247 500 281
rect 626 255 660 349
rect -660 187 -626 221
rect -660 119 -626 153
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect -660 -153 -626 -119
rect -660 -221 -626 -187
rect -546 187 -512 204
rect -546 119 -512 127
rect -546 51 -512 55
rect -546 -55 -512 -51
rect -546 -127 -512 -119
rect -546 -204 -512 -187
rect 512 187 546 204
rect 512 119 546 127
rect 512 51 546 55
rect 512 -55 546 -51
rect 512 -127 546 -119
rect 512 -204 546 -187
rect 626 187 660 221
rect 626 119 660 153
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect 626 -153 660 -119
rect 626 -221 660 -187
rect -660 -349 -626 -255
rect -500 -281 -459 -247
rect -415 -281 -391 -247
rect -343 -281 -323 -247
rect -271 -281 -255 -247
rect -199 -281 -187 -247
rect -127 -281 -119 -247
rect -55 -281 -51 -247
rect 51 -281 55 -247
rect 119 -281 127 -247
rect 187 -281 199 -247
rect 255 -281 271 -247
rect 323 -281 343 -247
rect 391 -281 415 -247
rect 459 -281 500 -247
rect 626 -349 660 -255
rect -660 -383 -561 -349
rect -527 -383 -493 -349
rect -459 -383 -425 -349
rect -391 -383 -357 -349
rect -323 -383 -289 -349
rect -255 -383 -221 -349
rect -187 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 187 -349
rect 221 -383 255 -349
rect 289 -383 323 -349
rect 357 -383 391 -349
rect 425 -383 459 -349
rect 493 -383 527 -349
rect 561 -383 660 -349
<< viali >>
rect -449 247 -425 281
rect -425 247 -415 281
rect -377 247 -357 281
rect -357 247 -343 281
rect -305 247 -289 281
rect -289 247 -271 281
rect -233 247 -221 281
rect -221 247 -199 281
rect -161 247 -153 281
rect -153 247 -127 281
rect -89 247 -85 281
rect -85 247 -55 281
rect -17 247 17 281
rect 55 247 85 281
rect 85 247 89 281
rect 127 247 153 281
rect 153 247 161 281
rect 199 247 221 281
rect 221 247 233 281
rect 271 247 289 281
rect 289 247 305 281
rect 343 247 357 281
rect 357 247 377 281
rect 415 247 425 281
rect 425 247 449 281
rect -546 153 -512 161
rect -546 127 -512 153
rect -546 85 -512 89
rect -546 55 -512 85
rect -546 -17 -512 17
rect -546 -85 -512 -55
rect -546 -89 -512 -85
rect -546 -153 -512 -127
rect -546 -161 -512 -153
rect 512 153 546 161
rect 512 127 546 153
rect 512 85 546 89
rect 512 55 546 85
rect 512 -17 546 17
rect 512 -85 546 -55
rect 512 -89 546 -85
rect 512 -153 546 -127
rect 512 -161 546 -153
rect -449 -281 -425 -247
rect -425 -281 -415 -247
rect -377 -281 -357 -247
rect -357 -281 -343 -247
rect -305 -281 -289 -247
rect -289 -281 -271 -247
rect -233 -281 -221 -247
rect -221 -281 -199 -247
rect -161 -281 -153 -247
rect -153 -281 -127 -247
rect -89 -281 -85 -247
rect -85 -281 -55 -247
rect -17 -281 17 -247
rect 55 -281 85 -247
rect 85 -281 89 -247
rect 127 -281 153 -247
rect 153 -281 161 -247
rect 199 -281 221 -247
rect 221 -281 233 -247
rect 271 -281 289 -247
rect 289 -281 305 -247
rect 343 -281 357 -247
rect 357 -281 377 -247
rect 415 -281 425 -247
rect 425 -281 449 -247
<< metal1 >>
rect -496 281 496 287
rect -496 247 -449 281
rect -415 247 -377 281
rect -343 247 -305 281
rect -271 247 -233 281
rect -199 247 -161 281
rect -127 247 -89 281
rect -55 247 -17 281
rect 17 247 55 281
rect 89 247 127 281
rect 161 247 199 281
rect 233 247 271 281
rect 305 247 343 281
rect 377 247 415 281
rect 449 247 496 281
rect -496 241 496 247
rect -552 161 -506 200
rect -552 127 -546 161
rect -512 127 -506 161
rect -552 89 -506 127
rect -552 55 -546 89
rect -512 55 -506 89
rect -552 17 -506 55
rect -552 -17 -546 17
rect -512 -17 -506 17
rect -552 -55 -506 -17
rect -552 -89 -546 -55
rect -512 -89 -506 -55
rect -552 -127 -506 -89
rect -552 -161 -546 -127
rect -512 -161 -506 -127
rect -552 -200 -506 -161
rect 506 161 552 200
rect 506 127 512 161
rect 546 127 552 161
rect 506 89 552 127
rect 506 55 512 89
rect 546 55 552 89
rect 506 17 552 55
rect 506 -17 512 17
rect 546 -17 552 17
rect 506 -55 552 -17
rect 506 -89 512 -55
rect 546 -89 552 -55
rect 506 -127 552 -89
rect 506 -161 512 -127
rect 546 -161 552 -127
rect 506 -200 552 -161
rect -496 -247 496 -241
rect -496 -281 -449 -247
rect -415 -281 -377 -247
rect -343 -281 -305 -247
rect -271 -281 -233 -247
rect -199 -281 -161 -247
rect -127 -281 -89 -247
rect -55 -281 -17 -247
rect 17 -281 55 -247
rect 89 -281 127 -247
rect 161 -281 199 -247
rect 233 -281 271 -247
rect 305 -281 343 -247
rect 377 -281 415 -247
rect 449 -281 496 -247
rect -496 -287 496 -281
<< properties >>
string FIXED_BBOX -643 -366 643 366
<< end >>
