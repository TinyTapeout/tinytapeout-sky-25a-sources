magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< error_p >>
rect -77 372 -19 378
rect 115 372 173 378
rect -77 338 -65 372
rect 115 338 127 372
rect -77 332 -19 338
rect 115 332 173 338
rect -173 -338 -115 -332
rect 19 -338 77 -332
rect -173 -372 -161 -338
rect 19 -372 31 -338
rect -173 -378 -115 -372
rect 19 -378 77 -372
<< pwell >>
rect -349 -500 349 500
<< nmos >>
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
<< ndiff >>
rect -221 255 -159 300
rect -221 221 -209 255
rect -175 221 -159 255
rect -221 187 -159 221
rect -221 153 -209 187
rect -175 153 -159 187
rect -221 119 -159 153
rect -221 85 -209 119
rect -175 85 -159 119
rect -221 51 -159 85
rect -221 17 -209 51
rect -175 17 -159 51
rect -221 -17 -159 17
rect -221 -51 -209 -17
rect -175 -51 -159 -17
rect -221 -85 -159 -51
rect -221 -119 -209 -85
rect -175 -119 -159 -85
rect -221 -153 -159 -119
rect -221 -187 -209 -153
rect -175 -187 -159 -153
rect -221 -221 -159 -187
rect -221 -255 -209 -221
rect -175 -255 -159 -221
rect -221 -300 -159 -255
rect -129 255 -63 300
rect -129 221 -113 255
rect -79 221 -63 255
rect -129 187 -63 221
rect -129 153 -113 187
rect -79 153 -63 187
rect -129 119 -63 153
rect -129 85 -113 119
rect -79 85 -63 119
rect -129 51 -63 85
rect -129 17 -113 51
rect -79 17 -63 51
rect -129 -17 -63 17
rect -129 -51 -113 -17
rect -79 -51 -63 -17
rect -129 -85 -63 -51
rect -129 -119 -113 -85
rect -79 -119 -63 -85
rect -129 -153 -63 -119
rect -129 -187 -113 -153
rect -79 -187 -63 -153
rect -129 -221 -63 -187
rect -129 -255 -113 -221
rect -79 -255 -63 -221
rect -129 -300 -63 -255
rect -33 255 33 300
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -300 33 -255
rect 63 255 129 300
rect 63 221 79 255
rect 113 221 129 255
rect 63 187 129 221
rect 63 153 79 187
rect 113 153 129 187
rect 63 119 129 153
rect 63 85 79 119
rect 113 85 129 119
rect 63 51 129 85
rect 63 17 79 51
rect 113 17 129 51
rect 63 -17 129 17
rect 63 -51 79 -17
rect 113 -51 129 -17
rect 63 -85 129 -51
rect 63 -119 79 -85
rect 113 -119 129 -85
rect 63 -153 129 -119
rect 63 -187 79 -153
rect 113 -187 129 -153
rect 63 -221 129 -187
rect 63 -255 79 -221
rect 113 -255 129 -221
rect 63 -300 129 -255
rect 159 255 221 300
rect 159 221 175 255
rect 209 221 221 255
rect 159 187 221 221
rect 159 153 175 187
rect 209 153 221 187
rect 159 119 221 153
rect 159 85 175 119
rect 209 85 221 119
rect 159 51 221 85
rect 159 17 175 51
rect 209 17 221 51
rect 159 -17 221 17
rect 159 -51 175 -17
rect 209 -51 221 -17
rect 159 -85 221 -51
rect 159 -119 175 -85
rect 209 -119 221 -85
rect 159 -153 221 -119
rect 159 -187 175 -153
rect 209 -187 221 -153
rect 159 -221 221 -187
rect 159 -255 175 -221
rect 209 -255 221 -221
rect 159 -300 221 -255
<< ndiffc >>
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
<< psubdiff >>
rect -323 440 -221 474
rect -187 440 -153 474
rect -119 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 119 474
rect 153 440 187 474
rect 221 440 323 474
rect -323 357 -289 440
rect -323 289 -289 323
rect 289 357 323 440
rect -323 221 -289 255
rect -323 153 -289 187
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect -323 -187 -289 -153
rect -323 -255 -289 -221
rect -323 -323 -289 -289
rect 289 289 323 323
rect 289 221 323 255
rect 289 153 323 187
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect 289 -119 323 -85
rect 289 -187 323 -153
rect 289 -255 323 -221
rect -323 -440 -289 -357
rect 289 -323 323 -289
rect 289 -440 323 -357
rect -323 -474 -221 -440
rect -187 -474 -153 -440
rect -119 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 119 -440
rect 153 -474 187 -440
rect 221 -474 323 -440
<< psubdiffcont >>
rect -221 440 -187 474
rect -153 440 -119 474
rect -85 440 -51 474
rect -17 440 17 474
rect 51 440 85 474
rect 119 440 153 474
rect 187 440 221 474
rect -323 323 -289 357
rect 289 323 323 357
rect -323 255 -289 289
rect -323 187 -289 221
rect -323 119 -289 153
rect -323 51 -289 85
rect -323 -17 -289 17
rect -323 -85 -289 -51
rect -323 -153 -289 -119
rect -323 -221 -289 -187
rect -323 -289 -289 -255
rect 289 255 323 289
rect 289 187 323 221
rect 289 119 323 153
rect 289 51 323 85
rect 289 -17 323 17
rect 289 -85 323 -51
rect 289 -153 323 -119
rect 289 -221 323 -187
rect 289 -289 323 -255
rect -323 -357 -289 -323
rect 289 -357 323 -323
rect -221 -474 -187 -440
rect -153 -474 -119 -440
rect -85 -474 -51 -440
rect -17 -474 17 -440
rect 51 -474 85 -440
rect 119 -474 153 -440
rect 187 -474 221 -440
<< poly >>
rect -81 372 -15 388
rect -81 338 -65 372
rect -31 338 -15 372
rect -159 300 -129 326
rect -81 322 -15 338
rect 111 372 177 388
rect 111 338 127 372
rect 161 338 177 372
rect -63 300 -33 322
rect 33 300 63 326
rect 111 322 177 338
rect 129 300 159 322
rect -159 -322 -129 -300
rect -177 -338 -111 -322
rect -63 -326 -33 -300
rect 33 -322 63 -300
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect -177 -388 -111 -372
rect 15 -338 81 -322
rect 129 -326 159 -300
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 15 -388 81 -372
<< polycont >>
rect -65 338 -31 372
rect 127 338 161 372
rect -161 -372 -127 -338
rect 31 -372 65 -338
<< locali >>
rect -323 440 -221 474
rect -187 440 -153 474
rect -119 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 119 474
rect 153 440 187 474
rect 221 440 323 474
rect -323 357 -289 440
rect -81 338 -65 372
rect -31 338 -15 372
rect 111 338 127 372
rect 161 338 177 372
rect 289 357 323 440
rect -323 289 -289 323
rect -323 221 -289 255
rect -323 153 -289 187
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect -323 -187 -289 -153
rect -323 -255 -289 -221
rect -323 -323 -289 -289
rect -209 269 -175 304
rect -209 197 -175 221
rect -209 125 -175 153
rect -209 53 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -53
rect -209 -153 -175 -125
rect -209 -221 -175 -197
rect -209 -304 -175 -269
rect -113 269 -79 304
rect -113 197 -79 221
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -221 -79 -197
rect -113 -304 -79 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 79 269 113 304
rect 79 197 113 221
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -221 113 -197
rect 79 -304 113 -269
rect 175 269 209 304
rect 175 197 209 221
rect 175 125 209 153
rect 175 53 209 85
rect 175 -17 209 17
rect 175 -85 209 -53
rect 175 -153 209 -125
rect 175 -221 209 -197
rect 175 -304 209 -269
rect 289 289 323 323
rect 289 221 323 255
rect 289 153 323 187
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect 289 -119 323 -85
rect 289 -187 323 -153
rect 289 -255 323 -221
rect 289 -323 323 -289
rect -323 -440 -289 -357
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 289 -440 323 -357
rect -323 -474 -221 -440
rect -187 -474 -153 -440
rect -119 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 119 -440
rect 153 -474 187 -440
rect 221 -474 323 -440
<< viali >>
rect -65 338 -31 372
rect 127 338 161 372
rect -209 255 -175 269
rect -209 235 -175 255
rect -209 187 -175 197
rect -209 163 -175 187
rect -209 119 -175 125
rect -209 91 -175 119
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -209 -119 -175 -91
rect -209 -125 -175 -119
rect -209 -187 -175 -163
rect -209 -197 -175 -187
rect -209 -255 -175 -235
rect -209 -269 -175 -255
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 175 255 209 269
rect 175 235 209 255
rect 175 187 209 197
rect 175 163 209 187
rect 175 119 209 125
rect 175 91 209 119
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 175 -119 209 -91
rect 175 -125 209 -119
rect 175 -187 209 -163
rect 175 -197 209 -187
rect 175 -255 209 -235
rect 175 -269 209 -255
rect -161 -372 -127 -338
rect 31 -372 65 -338
<< metal1 >>
rect -77 372 -19 378
rect -77 338 -65 372
rect -31 338 -19 372
rect -77 332 -19 338
rect 115 372 173 378
rect 115 338 127 372
rect 161 338 173 372
rect 115 332 173 338
rect -215 269 -169 300
rect -215 235 -209 269
rect -175 235 -169 269
rect -215 197 -169 235
rect -215 163 -209 197
rect -175 163 -169 197
rect -215 125 -169 163
rect -215 91 -209 125
rect -175 91 -169 125
rect -215 53 -169 91
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -91 -169 -53
rect -215 -125 -209 -91
rect -175 -125 -169 -91
rect -215 -163 -169 -125
rect -215 -197 -209 -163
rect -175 -197 -169 -163
rect -215 -235 -169 -197
rect -215 -269 -209 -235
rect -175 -269 -169 -235
rect -215 -300 -169 -269
rect -119 269 -73 300
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -300 -73 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 73 269 119 300
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -300 119 -269
rect 169 269 215 300
rect 169 235 175 269
rect 209 235 215 269
rect 169 197 215 235
rect 169 163 175 197
rect 209 163 215 197
rect 169 125 215 163
rect 169 91 175 125
rect 209 91 215 125
rect 169 53 215 91
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -91 215 -53
rect 169 -125 175 -91
rect 209 -125 215 -91
rect 169 -163 215 -125
rect 169 -197 175 -163
rect 209 -197 215 -163
rect 169 -235 215 -197
rect 169 -269 175 -235
rect 209 -269 215 -235
rect 169 -300 215 -269
rect -173 -338 -115 -332
rect -173 -372 -161 -338
rect -127 -372 -115 -338
rect -173 -378 -115 -372
rect 19 -338 77 -332
rect 19 -372 31 -338
rect 65 -372 77 -338
rect 19 -378 77 -372
<< properties >>
string FIXED_BBOX -306 -457 306 457
<< end >>
