magic
tech sky130A
magscale 1 1
timestamp 1740610800
<< checkpaint >>
rect 0 0 1664 1280
use JNWATR_NCH_12CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 832 240
use JNWATR_NCH_12C1F2 xa2 
transform 1 0 0 0 1 240
box 0 240 832 640
use JNWATR_NCH_12C5F0 xa3 
transform 1 0 0 0 1 640
box 0 640 832 1040
use JNWATR_NCH_12CTAPTOP xa4 
transform 1 0 0 0 1 1040
box 0 1040 832 1280
use JNWATR_NCH_12CTAPBOT xb1 
transform 1 0 832 0 1 0
box 832 0 1664 240
use JNWATR_NCH_12C1F2 xb2 
transform 1 0 832 0 1 240
box 832 240 1664 640
use JNWATR_NCH_12C5F0 xb3 
transform 1 0 832 0 1 640
box 832 640 1664 1040
use JNWATR_NCH_12CTAPTOP xb4 
transform 1 0 832 0 1 1040
box 832 1040 1664 1280
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1664 1280
<< end >>
