magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -189 1200 189 1286
rect -189 -1200 -103 1200
rect 103 -1200 189 1200
rect -189 -1286 189 -1200
<< psubdiff >>
rect -163 1226 -51 1260
rect -17 1226 17 1260
rect 51 1226 163 1260
rect -163 1139 -129 1226
rect 129 1139 163 1226
rect -163 1071 -129 1105
rect -163 1003 -129 1037
rect -163 935 -129 969
rect -163 867 -129 901
rect -163 799 -129 833
rect -163 731 -129 765
rect -163 663 -129 697
rect -163 595 -129 629
rect -163 527 -129 561
rect -163 459 -129 493
rect -163 391 -129 425
rect -163 323 -129 357
rect -163 255 -129 289
rect -163 187 -129 221
rect -163 119 -129 153
rect -163 51 -129 85
rect -163 -17 -129 17
rect -163 -85 -129 -51
rect -163 -153 -129 -119
rect -163 -221 -129 -187
rect -163 -289 -129 -255
rect -163 -357 -129 -323
rect -163 -425 -129 -391
rect -163 -493 -129 -459
rect -163 -561 -129 -527
rect -163 -629 -129 -595
rect -163 -697 -129 -663
rect -163 -765 -129 -731
rect -163 -833 -129 -799
rect -163 -901 -129 -867
rect -163 -969 -129 -935
rect -163 -1037 -129 -1003
rect -163 -1105 -129 -1071
rect 129 1071 163 1105
rect 129 1003 163 1037
rect 129 935 163 969
rect 129 867 163 901
rect 129 799 163 833
rect 129 731 163 765
rect 129 663 163 697
rect 129 595 163 629
rect 129 527 163 561
rect 129 459 163 493
rect 129 391 163 425
rect 129 323 163 357
rect 129 255 163 289
rect 129 187 163 221
rect 129 119 163 153
rect 129 51 163 85
rect 129 -17 163 17
rect 129 -85 163 -51
rect 129 -153 163 -119
rect 129 -221 163 -187
rect 129 -289 163 -255
rect 129 -357 163 -323
rect 129 -425 163 -391
rect 129 -493 163 -459
rect 129 -561 163 -527
rect 129 -629 163 -595
rect 129 -697 163 -663
rect 129 -765 163 -731
rect 129 -833 163 -799
rect 129 -901 163 -867
rect 129 -969 163 -935
rect 129 -1037 163 -1003
rect 129 -1105 163 -1071
rect -163 -1226 -129 -1139
rect 129 -1226 163 -1139
rect -163 -1260 -51 -1226
rect -17 -1260 17 -1226
rect 51 -1260 163 -1226
<< psubdiffcont >>
rect -51 1226 -17 1260
rect 17 1226 51 1260
rect -163 1105 -129 1139
rect -163 1037 -129 1071
rect -163 969 -129 1003
rect -163 901 -129 935
rect -163 833 -129 867
rect -163 765 -129 799
rect -163 697 -129 731
rect -163 629 -129 663
rect -163 561 -129 595
rect -163 493 -129 527
rect -163 425 -129 459
rect -163 357 -129 391
rect -163 289 -129 323
rect -163 221 -129 255
rect -163 153 -129 187
rect -163 85 -129 119
rect -163 17 -129 51
rect -163 -51 -129 -17
rect -163 -119 -129 -85
rect -163 -187 -129 -153
rect -163 -255 -129 -221
rect -163 -323 -129 -289
rect -163 -391 -129 -357
rect -163 -459 -129 -425
rect -163 -527 -129 -493
rect -163 -595 -129 -561
rect -163 -663 -129 -629
rect -163 -731 -129 -697
rect -163 -799 -129 -765
rect -163 -867 -129 -833
rect -163 -935 -129 -901
rect -163 -1003 -129 -969
rect -163 -1071 -129 -1037
rect -163 -1139 -129 -1105
rect 129 1105 163 1139
rect 129 1037 163 1071
rect 129 969 163 1003
rect 129 901 163 935
rect 129 833 163 867
rect 129 765 163 799
rect 129 697 163 731
rect 129 629 163 663
rect 129 561 163 595
rect 129 493 163 527
rect 129 425 163 459
rect 129 357 163 391
rect 129 289 163 323
rect 129 221 163 255
rect 129 153 163 187
rect 129 85 163 119
rect 129 17 163 51
rect 129 -51 163 -17
rect 129 -119 163 -85
rect 129 -187 163 -153
rect 129 -255 163 -221
rect 129 -323 163 -289
rect 129 -391 163 -357
rect 129 -459 163 -425
rect 129 -527 163 -493
rect 129 -595 163 -561
rect 129 -663 163 -629
rect 129 -731 163 -697
rect 129 -799 163 -765
rect 129 -867 163 -833
rect 129 -935 163 -901
rect 129 -1003 163 -969
rect 129 -1071 163 -1037
rect 129 -1139 163 -1105
rect -51 -1260 -17 -1226
rect 17 -1260 51 -1226
<< poly >>
rect -33 1114 33 1130
rect -33 1080 -17 1114
rect 17 1080 33 1114
rect -33 700 33 1080
rect -33 -1080 33 -700
rect -33 -1114 -17 -1080
rect 17 -1114 33 -1080
rect -33 -1130 33 -1114
<< polycont >>
rect -17 1080 17 1114
rect -17 -1114 17 -1080
<< npolyres >>
rect -33 -700 33 700
<< locali >>
rect -163 1226 -51 1260
rect -17 1226 17 1260
rect 51 1226 163 1260
rect -163 1139 -129 1226
rect 129 1139 163 1226
rect -163 1071 -129 1105
rect -33 1080 -17 1114
rect 17 1080 33 1114
rect -163 1003 -129 1037
rect -163 935 -129 969
rect -163 867 -129 901
rect -163 799 -129 833
rect -163 731 -129 765
rect -17 1040 17 1078
rect -17 968 17 1006
rect -17 896 17 934
rect -17 824 17 862
rect -17 752 17 790
rect -17 717 17 718
rect 129 1071 163 1105
rect 129 1003 163 1037
rect 129 935 163 969
rect 129 867 163 901
rect 129 799 163 833
rect 129 731 163 765
rect -163 663 -129 697
rect -163 595 -129 629
rect -163 527 -129 561
rect -163 459 -129 493
rect -163 391 -129 425
rect -163 323 -129 357
rect -163 255 -129 289
rect -163 187 -129 221
rect -163 119 -129 153
rect -163 51 -129 85
rect -163 -17 -129 17
rect -163 -85 -129 -51
rect -163 -153 -129 -119
rect -163 -221 -129 -187
rect -163 -289 -129 -255
rect -163 -357 -129 -323
rect -163 -425 -129 -391
rect -163 -493 -129 -459
rect -163 -561 -129 -527
rect -163 -629 -129 -595
rect -163 -697 -129 -663
rect 129 663 163 697
rect 129 595 163 629
rect 129 527 163 561
rect 129 459 163 493
rect 129 391 163 425
rect 129 323 163 357
rect 129 255 163 289
rect 129 187 163 221
rect 129 119 163 153
rect 129 51 163 85
rect 129 -17 163 17
rect 129 -85 163 -51
rect 129 -153 163 -119
rect 129 -221 163 -187
rect 129 -289 163 -255
rect 129 -357 163 -323
rect 129 -425 163 -391
rect 129 -493 163 -459
rect 129 -561 163 -527
rect 129 -629 163 -595
rect 129 -697 163 -663
rect -163 -765 -129 -731
rect -163 -833 -129 -799
rect -163 -901 -129 -867
rect -163 -969 -129 -935
rect -163 -1037 -129 -1003
rect -163 -1105 -129 -1071
rect -17 -719 17 -717
rect -17 -791 17 -753
rect -17 -863 17 -825
rect -17 -935 17 -897
rect -17 -1007 17 -969
rect -17 -1079 17 -1041
rect 129 -765 163 -731
rect 129 -833 163 -799
rect 129 -901 163 -867
rect 129 -969 163 -935
rect 129 -1037 163 -1003
rect -33 -1114 -17 -1080
rect 17 -1114 33 -1080
rect 129 -1105 163 -1071
rect -163 -1226 -129 -1139
rect 129 -1226 163 -1139
rect -163 -1260 -51 -1226
rect -17 -1260 17 -1226
rect 51 -1260 163 -1226
<< viali >>
rect -17 1080 17 1112
rect -17 1078 17 1080
rect -17 1006 17 1040
rect -17 934 17 968
rect -17 862 17 896
rect -17 790 17 824
rect -17 718 17 752
rect -17 -753 17 -719
rect -17 -825 17 -791
rect -17 -897 17 -863
rect -17 -969 17 -935
rect -17 -1041 17 -1007
rect -17 -1080 17 -1079
rect -17 -1113 17 -1080
<< metal1 >>
rect -23 1112 23 1126
rect -23 1078 -17 1112
rect 17 1078 23 1112
rect -23 1040 23 1078
rect -23 1006 -17 1040
rect 17 1006 23 1040
rect -23 968 23 1006
rect -23 934 -17 968
rect 17 934 23 968
rect -23 896 23 934
rect -23 862 -17 896
rect 17 862 23 896
rect -23 824 23 862
rect -23 790 -17 824
rect 17 790 23 824
rect -23 752 23 790
rect -23 718 -17 752
rect 17 718 23 752
rect -23 705 23 718
rect -23 -719 23 -705
rect -23 -753 -17 -719
rect 17 -753 23 -719
rect -23 -791 23 -753
rect -23 -825 -17 -791
rect 17 -825 23 -791
rect -23 -863 23 -825
rect -23 -897 -17 -863
rect 17 -897 23 -863
rect -23 -935 23 -897
rect -23 -969 -17 -935
rect 17 -969 23 -935
rect -23 -1007 23 -969
rect -23 -1041 -17 -1007
rect 17 -1041 23 -1007
rect -23 -1079 23 -1041
rect -23 -1113 -17 -1079
rect 17 -1113 23 -1079
rect -23 -1126 23 -1113
<< properties >>
string FIXED_BBOX -146 -1243 146 1243
<< end >>
