magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< pwell >>
rect -225 676 225 762
rect -225 -676 -139 676
rect 139 -676 225 676
rect -225 -762 225 -676
<< psubdiff >>
rect -199 702 -85 736
rect -51 702 -17 736
rect 17 702 51 736
rect 85 702 199 736
rect -199 629 -165 702
rect 165 629 199 702
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect -199 -702 -165 -629
rect 165 -702 199 -629
rect -199 -736 -85 -702
rect -51 -736 -17 -702
rect 17 -736 51 -702
rect 85 -736 199 -702
<< psubdiffcont >>
rect -85 702 -51 736
rect -17 702 17 736
rect 51 702 85 736
rect -199 595 -165 629
rect -199 527 -165 561
rect -199 459 -165 493
rect -199 391 -165 425
rect -199 323 -165 357
rect -199 255 -165 289
rect -199 187 -165 221
rect -199 119 -165 153
rect -199 51 -165 85
rect -199 -17 -165 17
rect -199 -85 -165 -51
rect -199 -153 -165 -119
rect -199 -221 -165 -187
rect -199 -289 -165 -255
rect -199 -357 -165 -323
rect -199 -425 -165 -391
rect -199 -493 -165 -459
rect -199 -561 -165 -527
rect -199 -629 -165 -595
rect 165 595 199 629
rect 165 527 199 561
rect 165 459 199 493
rect 165 391 199 425
rect 165 323 199 357
rect 165 255 199 289
rect 165 187 199 221
rect 165 119 199 153
rect 165 51 199 85
rect 165 -17 199 17
rect 165 -85 199 -51
rect 165 -153 199 -119
rect 165 -221 199 -187
rect 165 -289 199 -255
rect 165 -357 199 -323
rect 165 -425 199 -391
rect 165 -493 199 -459
rect 165 -561 199 -527
rect 165 -629 199 -595
rect -85 -736 -51 -702
rect -17 -736 17 -702
rect 51 -736 85 -702
<< xpolycontact >>
rect -69 174 69 606
rect -69 -606 69 -174
<< ppolyres >>
rect -69 -174 69 174
<< locali >>
rect -199 702 -85 736
rect -51 702 -17 736
rect 17 702 51 736
rect 85 702 199 736
rect -199 629 -165 702
rect 165 629 199 702
rect -199 561 -165 595
rect -199 493 -165 527
rect -199 425 -165 459
rect -199 357 -165 391
rect -199 289 -165 323
rect -199 221 -165 255
rect -199 153 -165 187
rect 165 561 199 595
rect 165 493 199 527
rect 165 425 199 459
rect 165 357 199 391
rect 165 289 199 323
rect 165 221 199 255
rect -199 85 -165 119
rect -199 17 -165 51
rect -199 -51 -165 -17
rect -199 -119 -165 -85
rect -199 -187 -165 -153
rect 165 153 199 187
rect 165 85 199 119
rect 165 17 199 51
rect 165 -51 199 -17
rect 165 -119 199 -85
rect -199 -255 -165 -221
rect -199 -323 -165 -289
rect -199 -391 -165 -357
rect -199 -459 -165 -425
rect -199 -527 -165 -493
rect -199 -595 -165 -561
rect 165 -187 199 -153
rect 165 -255 199 -221
rect 165 -323 199 -289
rect 165 -391 199 -357
rect 165 -459 199 -425
rect 165 -527 199 -493
rect 165 -595 199 -561
rect -199 -702 -165 -629
rect 165 -702 199 -629
rect -199 -736 -85 -702
rect -51 -736 -17 -702
rect 17 -736 51 -702
rect 85 -736 199 -702
<< viali >>
rect -53 192 53 586
<< metal1 >>
rect -59 586 59 600
rect -59 192 -53 586
rect 53 192 59 586
rect -59 179 59 192
rect -59 -600 59 -179
<< properties >>
string FIXED_BBOX -182 -719 182 719
<< end >>
