magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< metal3 >>
rect -3186 2992 3186 3040
rect -3186 2928 3102 2992
rect 3166 2928 3186 2992
rect -3186 2912 3186 2928
rect -3186 2848 3102 2912
rect 3166 2848 3186 2912
rect -3186 2832 3186 2848
rect -3186 2768 3102 2832
rect 3166 2768 3186 2832
rect -3186 2752 3186 2768
rect -3186 2688 3102 2752
rect 3166 2688 3186 2752
rect -3186 2672 3186 2688
rect -3186 2608 3102 2672
rect 3166 2608 3186 2672
rect -3186 2592 3186 2608
rect -3186 2528 3102 2592
rect 3166 2528 3186 2592
rect -3186 2512 3186 2528
rect -3186 2448 3102 2512
rect 3166 2448 3186 2512
rect -3186 2432 3186 2448
rect -3186 2368 3102 2432
rect 3166 2368 3186 2432
rect -3186 2352 3186 2368
rect -3186 2288 3102 2352
rect 3166 2288 3186 2352
rect -3186 2272 3186 2288
rect -3186 2208 3102 2272
rect 3166 2208 3186 2272
rect -3186 2192 3186 2208
rect -3186 2128 3102 2192
rect 3166 2128 3186 2192
rect -3186 2112 3186 2128
rect -3186 2048 3102 2112
rect 3166 2048 3186 2112
rect -3186 2032 3186 2048
rect -3186 1968 3102 2032
rect 3166 1968 3186 2032
rect -3186 1952 3186 1968
rect -3186 1888 3102 1952
rect 3166 1888 3186 1952
rect -3186 1872 3186 1888
rect -3186 1808 3102 1872
rect 3166 1808 3186 1872
rect -3186 1792 3186 1808
rect -3186 1728 3102 1792
rect 3166 1728 3186 1792
rect -3186 1712 3186 1728
rect -3186 1648 3102 1712
rect 3166 1648 3186 1712
rect -3186 1632 3186 1648
rect -3186 1568 3102 1632
rect 3166 1568 3186 1632
rect -3186 1552 3186 1568
rect -3186 1488 3102 1552
rect 3166 1488 3186 1552
rect -3186 1472 3186 1488
rect -3186 1408 3102 1472
rect 3166 1408 3186 1472
rect -3186 1392 3186 1408
rect -3186 1328 3102 1392
rect 3166 1328 3186 1392
rect -3186 1312 3186 1328
rect -3186 1248 3102 1312
rect 3166 1248 3186 1312
rect -3186 1232 3186 1248
rect -3186 1168 3102 1232
rect 3166 1168 3186 1232
rect -3186 1152 3186 1168
rect -3186 1088 3102 1152
rect 3166 1088 3186 1152
rect -3186 1072 3186 1088
rect -3186 1008 3102 1072
rect 3166 1008 3186 1072
rect -3186 992 3186 1008
rect -3186 928 3102 992
rect 3166 928 3186 992
rect -3186 912 3186 928
rect -3186 848 3102 912
rect 3166 848 3186 912
rect -3186 832 3186 848
rect -3186 768 3102 832
rect 3166 768 3186 832
rect -3186 752 3186 768
rect -3186 688 3102 752
rect 3166 688 3186 752
rect -3186 672 3186 688
rect -3186 608 3102 672
rect 3166 608 3186 672
rect -3186 592 3186 608
rect -3186 528 3102 592
rect 3166 528 3186 592
rect -3186 512 3186 528
rect -3186 448 3102 512
rect 3166 448 3186 512
rect -3186 432 3186 448
rect -3186 368 3102 432
rect 3166 368 3186 432
rect -3186 352 3186 368
rect -3186 288 3102 352
rect 3166 288 3186 352
rect -3186 272 3186 288
rect -3186 208 3102 272
rect 3166 208 3186 272
rect -3186 192 3186 208
rect -3186 128 3102 192
rect 3166 128 3186 192
rect -3186 112 3186 128
rect -3186 48 3102 112
rect 3166 48 3186 112
rect -3186 32 3186 48
rect -3186 -32 3102 32
rect 3166 -32 3186 32
rect -3186 -48 3186 -32
rect -3186 -112 3102 -48
rect 3166 -112 3186 -48
rect -3186 -128 3186 -112
rect -3186 -192 3102 -128
rect 3166 -192 3186 -128
rect -3186 -208 3186 -192
rect -3186 -272 3102 -208
rect 3166 -272 3186 -208
rect -3186 -288 3186 -272
rect -3186 -352 3102 -288
rect 3166 -352 3186 -288
rect -3186 -368 3186 -352
rect -3186 -432 3102 -368
rect 3166 -432 3186 -368
rect -3186 -448 3186 -432
rect -3186 -512 3102 -448
rect 3166 -512 3186 -448
rect -3186 -528 3186 -512
rect -3186 -592 3102 -528
rect 3166 -592 3186 -528
rect -3186 -608 3186 -592
rect -3186 -672 3102 -608
rect 3166 -672 3186 -608
rect -3186 -688 3186 -672
rect -3186 -752 3102 -688
rect 3166 -752 3186 -688
rect -3186 -768 3186 -752
rect -3186 -832 3102 -768
rect 3166 -832 3186 -768
rect -3186 -848 3186 -832
rect -3186 -912 3102 -848
rect 3166 -912 3186 -848
rect -3186 -928 3186 -912
rect -3186 -992 3102 -928
rect 3166 -992 3186 -928
rect -3186 -1008 3186 -992
rect -3186 -1072 3102 -1008
rect 3166 -1072 3186 -1008
rect -3186 -1088 3186 -1072
rect -3186 -1152 3102 -1088
rect 3166 -1152 3186 -1088
rect -3186 -1168 3186 -1152
rect -3186 -1232 3102 -1168
rect 3166 -1232 3186 -1168
rect -3186 -1248 3186 -1232
rect -3186 -1312 3102 -1248
rect 3166 -1312 3186 -1248
rect -3186 -1328 3186 -1312
rect -3186 -1392 3102 -1328
rect 3166 -1392 3186 -1328
rect -3186 -1408 3186 -1392
rect -3186 -1472 3102 -1408
rect 3166 -1472 3186 -1408
rect -3186 -1488 3186 -1472
rect -3186 -1552 3102 -1488
rect 3166 -1552 3186 -1488
rect -3186 -1568 3186 -1552
rect -3186 -1632 3102 -1568
rect 3166 -1632 3186 -1568
rect -3186 -1648 3186 -1632
rect -3186 -1712 3102 -1648
rect 3166 -1712 3186 -1648
rect -3186 -1728 3186 -1712
rect -3186 -1792 3102 -1728
rect 3166 -1792 3186 -1728
rect -3186 -1808 3186 -1792
rect -3186 -1872 3102 -1808
rect 3166 -1872 3186 -1808
rect -3186 -1888 3186 -1872
rect -3186 -1952 3102 -1888
rect 3166 -1952 3186 -1888
rect -3186 -1968 3186 -1952
rect -3186 -2032 3102 -1968
rect 3166 -2032 3186 -1968
rect -3186 -2048 3186 -2032
rect -3186 -2112 3102 -2048
rect 3166 -2112 3186 -2048
rect -3186 -2128 3186 -2112
rect -3186 -2192 3102 -2128
rect 3166 -2192 3186 -2128
rect -3186 -2208 3186 -2192
rect -3186 -2272 3102 -2208
rect 3166 -2272 3186 -2208
rect -3186 -2288 3186 -2272
rect -3186 -2352 3102 -2288
rect 3166 -2352 3186 -2288
rect -3186 -2368 3186 -2352
rect -3186 -2432 3102 -2368
rect 3166 -2432 3186 -2368
rect -3186 -2448 3186 -2432
rect -3186 -2512 3102 -2448
rect 3166 -2512 3186 -2448
rect -3186 -2528 3186 -2512
rect -3186 -2592 3102 -2528
rect 3166 -2592 3186 -2528
rect -3186 -2608 3186 -2592
rect -3186 -2672 3102 -2608
rect 3166 -2672 3186 -2608
rect -3186 -2688 3186 -2672
rect -3186 -2752 3102 -2688
rect 3166 -2752 3186 -2688
rect -3186 -2768 3186 -2752
rect -3186 -2832 3102 -2768
rect 3166 -2832 3186 -2768
rect -3186 -2848 3186 -2832
rect -3186 -2912 3102 -2848
rect 3166 -2912 3186 -2848
rect -3186 -2928 3186 -2912
rect -3186 -2992 3102 -2928
rect 3166 -2992 3186 -2928
rect -3186 -3040 3186 -2992
<< via3 >>
rect 3102 2928 3166 2992
rect 3102 2848 3166 2912
rect 3102 2768 3166 2832
rect 3102 2688 3166 2752
rect 3102 2608 3166 2672
rect 3102 2528 3166 2592
rect 3102 2448 3166 2512
rect 3102 2368 3166 2432
rect 3102 2288 3166 2352
rect 3102 2208 3166 2272
rect 3102 2128 3166 2192
rect 3102 2048 3166 2112
rect 3102 1968 3166 2032
rect 3102 1888 3166 1952
rect 3102 1808 3166 1872
rect 3102 1728 3166 1792
rect 3102 1648 3166 1712
rect 3102 1568 3166 1632
rect 3102 1488 3166 1552
rect 3102 1408 3166 1472
rect 3102 1328 3166 1392
rect 3102 1248 3166 1312
rect 3102 1168 3166 1232
rect 3102 1088 3166 1152
rect 3102 1008 3166 1072
rect 3102 928 3166 992
rect 3102 848 3166 912
rect 3102 768 3166 832
rect 3102 688 3166 752
rect 3102 608 3166 672
rect 3102 528 3166 592
rect 3102 448 3166 512
rect 3102 368 3166 432
rect 3102 288 3166 352
rect 3102 208 3166 272
rect 3102 128 3166 192
rect 3102 48 3166 112
rect 3102 -32 3166 32
rect 3102 -112 3166 -48
rect 3102 -192 3166 -128
rect 3102 -272 3166 -208
rect 3102 -352 3166 -288
rect 3102 -432 3166 -368
rect 3102 -512 3166 -448
rect 3102 -592 3166 -528
rect 3102 -672 3166 -608
rect 3102 -752 3166 -688
rect 3102 -832 3166 -768
rect 3102 -912 3166 -848
rect 3102 -992 3166 -928
rect 3102 -1072 3166 -1008
rect 3102 -1152 3166 -1088
rect 3102 -1232 3166 -1168
rect 3102 -1312 3166 -1248
rect 3102 -1392 3166 -1328
rect 3102 -1472 3166 -1408
rect 3102 -1552 3166 -1488
rect 3102 -1632 3166 -1568
rect 3102 -1712 3166 -1648
rect 3102 -1792 3166 -1728
rect 3102 -1872 3166 -1808
rect 3102 -1952 3166 -1888
rect 3102 -2032 3166 -1968
rect 3102 -2112 3166 -2048
rect 3102 -2192 3166 -2128
rect 3102 -2272 3166 -2208
rect 3102 -2352 3166 -2288
rect 3102 -2432 3166 -2368
rect 3102 -2512 3166 -2448
rect 3102 -2592 3166 -2528
rect 3102 -2672 3166 -2608
rect 3102 -2752 3166 -2688
rect 3102 -2832 3166 -2768
rect 3102 -2912 3166 -2848
rect 3102 -2992 3166 -2928
<< mimcap >>
rect -3146 2952 2854 3000
rect -3146 -2952 -3098 2952
rect 2806 -2952 2854 2952
rect -3146 -3000 2854 -2952
<< mimcapcontact >>
rect -3098 -2952 2806 2952
<< metal4 >>
rect 3086 2992 3182 3028
rect -3107 2952 2815 2961
rect -3107 -2952 -3098 2952
rect 2806 -2952 2815 2952
rect -3107 -2961 2815 -2952
rect 3086 2928 3102 2992
rect 3166 2928 3182 2992
rect 3086 2912 3182 2928
rect 3086 2848 3102 2912
rect 3166 2848 3182 2912
rect 3086 2832 3182 2848
rect 3086 2768 3102 2832
rect 3166 2768 3182 2832
rect 3086 2752 3182 2768
rect 3086 2688 3102 2752
rect 3166 2688 3182 2752
rect 3086 2672 3182 2688
rect 3086 2608 3102 2672
rect 3166 2608 3182 2672
rect 3086 2592 3182 2608
rect 3086 2528 3102 2592
rect 3166 2528 3182 2592
rect 3086 2512 3182 2528
rect 3086 2448 3102 2512
rect 3166 2448 3182 2512
rect 3086 2432 3182 2448
rect 3086 2368 3102 2432
rect 3166 2368 3182 2432
rect 3086 2352 3182 2368
rect 3086 2288 3102 2352
rect 3166 2288 3182 2352
rect 3086 2272 3182 2288
rect 3086 2208 3102 2272
rect 3166 2208 3182 2272
rect 3086 2192 3182 2208
rect 3086 2128 3102 2192
rect 3166 2128 3182 2192
rect 3086 2112 3182 2128
rect 3086 2048 3102 2112
rect 3166 2048 3182 2112
rect 3086 2032 3182 2048
rect 3086 1968 3102 2032
rect 3166 1968 3182 2032
rect 3086 1952 3182 1968
rect 3086 1888 3102 1952
rect 3166 1888 3182 1952
rect 3086 1872 3182 1888
rect 3086 1808 3102 1872
rect 3166 1808 3182 1872
rect 3086 1792 3182 1808
rect 3086 1728 3102 1792
rect 3166 1728 3182 1792
rect 3086 1712 3182 1728
rect 3086 1648 3102 1712
rect 3166 1648 3182 1712
rect 3086 1632 3182 1648
rect 3086 1568 3102 1632
rect 3166 1568 3182 1632
rect 3086 1552 3182 1568
rect 3086 1488 3102 1552
rect 3166 1488 3182 1552
rect 3086 1472 3182 1488
rect 3086 1408 3102 1472
rect 3166 1408 3182 1472
rect 3086 1392 3182 1408
rect 3086 1328 3102 1392
rect 3166 1328 3182 1392
rect 3086 1312 3182 1328
rect 3086 1248 3102 1312
rect 3166 1248 3182 1312
rect 3086 1232 3182 1248
rect 3086 1168 3102 1232
rect 3166 1168 3182 1232
rect 3086 1152 3182 1168
rect 3086 1088 3102 1152
rect 3166 1088 3182 1152
rect 3086 1072 3182 1088
rect 3086 1008 3102 1072
rect 3166 1008 3182 1072
rect 3086 992 3182 1008
rect 3086 928 3102 992
rect 3166 928 3182 992
rect 3086 912 3182 928
rect 3086 848 3102 912
rect 3166 848 3182 912
rect 3086 832 3182 848
rect 3086 768 3102 832
rect 3166 768 3182 832
rect 3086 752 3182 768
rect 3086 688 3102 752
rect 3166 688 3182 752
rect 3086 672 3182 688
rect 3086 608 3102 672
rect 3166 608 3182 672
rect 3086 592 3182 608
rect 3086 528 3102 592
rect 3166 528 3182 592
rect 3086 512 3182 528
rect 3086 448 3102 512
rect 3166 448 3182 512
rect 3086 432 3182 448
rect 3086 368 3102 432
rect 3166 368 3182 432
rect 3086 352 3182 368
rect 3086 288 3102 352
rect 3166 288 3182 352
rect 3086 272 3182 288
rect 3086 208 3102 272
rect 3166 208 3182 272
rect 3086 192 3182 208
rect 3086 128 3102 192
rect 3166 128 3182 192
rect 3086 112 3182 128
rect 3086 48 3102 112
rect 3166 48 3182 112
rect 3086 32 3182 48
rect 3086 -32 3102 32
rect 3166 -32 3182 32
rect 3086 -48 3182 -32
rect 3086 -112 3102 -48
rect 3166 -112 3182 -48
rect 3086 -128 3182 -112
rect 3086 -192 3102 -128
rect 3166 -192 3182 -128
rect 3086 -208 3182 -192
rect 3086 -272 3102 -208
rect 3166 -272 3182 -208
rect 3086 -288 3182 -272
rect 3086 -352 3102 -288
rect 3166 -352 3182 -288
rect 3086 -368 3182 -352
rect 3086 -432 3102 -368
rect 3166 -432 3182 -368
rect 3086 -448 3182 -432
rect 3086 -512 3102 -448
rect 3166 -512 3182 -448
rect 3086 -528 3182 -512
rect 3086 -592 3102 -528
rect 3166 -592 3182 -528
rect 3086 -608 3182 -592
rect 3086 -672 3102 -608
rect 3166 -672 3182 -608
rect 3086 -688 3182 -672
rect 3086 -752 3102 -688
rect 3166 -752 3182 -688
rect 3086 -768 3182 -752
rect 3086 -832 3102 -768
rect 3166 -832 3182 -768
rect 3086 -848 3182 -832
rect 3086 -912 3102 -848
rect 3166 -912 3182 -848
rect 3086 -928 3182 -912
rect 3086 -992 3102 -928
rect 3166 -992 3182 -928
rect 3086 -1008 3182 -992
rect 3086 -1072 3102 -1008
rect 3166 -1072 3182 -1008
rect 3086 -1088 3182 -1072
rect 3086 -1152 3102 -1088
rect 3166 -1152 3182 -1088
rect 3086 -1168 3182 -1152
rect 3086 -1232 3102 -1168
rect 3166 -1232 3182 -1168
rect 3086 -1248 3182 -1232
rect 3086 -1312 3102 -1248
rect 3166 -1312 3182 -1248
rect 3086 -1328 3182 -1312
rect 3086 -1392 3102 -1328
rect 3166 -1392 3182 -1328
rect 3086 -1408 3182 -1392
rect 3086 -1472 3102 -1408
rect 3166 -1472 3182 -1408
rect 3086 -1488 3182 -1472
rect 3086 -1552 3102 -1488
rect 3166 -1552 3182 -1488
rect 3086 -1568 3182 -1552
rect 3086 -1632 3102 -1568
rect 3166 -1632 3182 -1568
rect 3086 -1648 3182 -1632
rect 3086 -1712 3102 -1648
rect 3166 -1712 3182 -1648
rect 3086 -1728 3182 -1712
rect 3086 -1792 3102 -1728
rect 3166 -1792 3182 -1728
rect 3086 -1808 3182 -1792
rect 3086 -1872 3102 -1808
rect 3166 -1872 3182 -1808
rect 3086 -1888 3182 -1872
rect 3086 -1952 3102 -1888
rect 3166 -1952 3182 -1888
rect 3086 -1968 3182 -1952
rect 3086 -2032 3102 -1968
rect 3166 -2032 3182 -1968
rect 3086 -2048 3182 -2032
rect 3086 -2112 3102 -2048
rect 3166 -2112 3182 -2048
rect 3086 -2128 3182 -2112
rect 3086 -2192 3102 -2128
rect 3166 -2192 3182 -2128
rect 3086 -2208 3182 -2192
rect 3086 -2272 3102 -2208
rect 3166 -2272 3182 -2208
rect 3086 -2288 3182 -2272
rect 3086 -2352 3102 -2288
rect 3166 -2352 3182 -2288
rect 3086 -2368 3182 -2352
rect 3086 -2432 3102 -2368
rect 3166 -2432 3182 -2368
rect 3086 -2448 3182 -2432
rect 3086 -2512 3102 -2448
rect 3166 -2512 3182 -2448
rect 3086 -2528 3182 -2512
rect 3086 -2592 3102 -2528
rect 3166 -2592 3182 -2528
rect 3086 -2608 3182 -2592
rect 3086 -2672 3102 -2608
rect 3166 -2672 3182 -2608
rect 3086 -2688 3182 -2672
rect 3086 -2752 3102 -2688
rect 3166 -2752 3182 -2688
rect 3086 -2768 3182 -2752
rect 3086 -2832 3102 -2768
rect 3166 -2832 3182 -2768
rect 3086 -2848 3182 -2832
rect 3086 -2912 3102 -2848
rect 3166 -2912 3182 -2848
rect 3086 -2928 3182 -2912
rect 3086 -2992 3102 -2928
rect 3166 -2992 3182 -2928
rect 3086 -3028 3182 -2992
<< properties >>
string FIXED_BBOX -3186 -3040 2894 3040
<< end >>
