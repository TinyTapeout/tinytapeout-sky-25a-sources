magic
tech sky130A
magscale 1 2
timestamp 1756992108
<< nwell >>
rect -296 -319 296 319
<< pmos >>
rect -100 -100 100 100
<< pdiff >>
rect -158 85 -100 100
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -100 -100 -85
rect 100 85 158 100
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -100 158 -85
<< pdiffc >>
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
<< nsubdiff >>
rect -260 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 260 283
rect -260 187 -226 249
rect -260 119 -226 153
rect 226 187 260 249
rect 226 119 260 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect -260 -153 -226 -119
rect -260 -249 -226 -187
rect 226 -153 260 -119
rect 226 -249 260 -187
rect -260 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 260 -249
<< nsubdiffcont >>
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect -260 153 -226 187
rect -260 85 -226 119
rect 226 153 260 187
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect -260 -187 -226 -153
rect 226 -119 260 -85
rect 226 -187 260 -153
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
<< poly >>
rect -100 181 100 197
rect -100 147 -51 181
rect -17 147 17 181
rect 51 147 100 181
rect -100 100 100 147
rect -100 -147 100 -100
rect -100 -181 -51 -147
rect -17 -181 17 -147
rect 51 -181 100 -147
rect -100 -197 100 -181
<< polycont >>
rect -51 147 -17 181
rect 17 147 51 181
rect -51 -181 -17 -147
rect 17 -181 51 -147
<< locali >>
rect -260 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 260 283
rect -260 187 -226 249
rect 226 187 260 249
rect -260 119 -226 153
rect -100 147 -53 181
rect -17 147 17 181
rect 53 147 100 181
rect 226 119 260 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -146 85 -112 104
rect -146 17 -112 19
rect -146 -19 -112 -17
rect -146 -104 -112 -85
rect 112 85 146 104
rect 112 17 146 19
rect 112 -19 146 -17
rect 112 -104 146 -85
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect -260 -153 -226 -119
rect -100 -181 -53 -147
rect -17 -181 17 -147
rect 53 -181 100 -147
rect 226 -153 260 -119
rect -260 -249 -226 -187
rect 226 -249 260 -187
rect -260 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 260 -249
<< viali >>
rect -53 147 -51 181
rect -51 147 -19 181
rect 19 147 51 181
rect 51 147 53 181
rect -146 51 -112 53
rect -146 19 -112 51
rect -146 -51 -112 -19
rect -146 -53 -112 -51
rect 112 51 146 53
rect 112 19 146 51
rect 112 -51 146 -19
rect 112 -53 146 -51
rect -53 -181 -51 -147
rect -51 -181 -19 -147
rect 19 -181 51 -147
rect 51 -181 53 -147
<< metal1 >>
rect -96 181 96 187
rect -96 147 -53 181
rect -19 147 19 181
rect 53 147 96 181
rect -96 141 96 147
rect -152 53 -106 100
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -100 -106 -53
rect 106 53 152 100
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -100 152 -53
rect -96 -147 96 -141
rect -96 -181 -53 -147
rect -19 -181 19 -147
rect 53 -181 96 -147
rect -96 -187 96 -181
<< properties >>
string FIXED_BBOX -243 -266 243 266
<< end >>
