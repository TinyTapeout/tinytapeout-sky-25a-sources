// Generated from: 20250609-230107_binTestAcc9746_seed1018940_epochs30_2x2560_b256_lr50_interconnect.pth

module net (
    input  wire [255:0] in,
    output wire [2559:0] out,
    output wire [1269:0] categories
);
    wire [2560:0] layer_0;

    // Layer 0 ============================================================
    assign layer_0[0] = ~(in[146] | in[150]); 
    assign layer_0[1] = in[228] | in[206]; 
    assign layer_0[2] = in[165] & ~in[250]; 
    assign layer_0[3] = in[107]; 
    assign layer_0[4] = in[105] & ~in[116]; 
    assign layer_0[5] = in[131] & ~in[215]; 
    assign layer_0[6] = in[57] & ~in[12]; 
    assign layer_0[7] = ~(in[85] ^ in[99]); 
    assign layer_0[8] = ~in[30]; 
    assign layer_0[9] = in[126]; 
    assign layer_0[10] = in[83] ^ in[53]; 
    assign layer_0[11] = in[119] ^ in[85]; 
    assign layer_0[12] = ~(in[137] ^ in[89]); 
    assign layer_0[13] = in[61] ^ in[108]; 
    assign layer_0[14] = in[210]; 
    assign layer_0[15] = ~in[26] | (in[26] & in[121]); 
    assign layer_0[16] = ~(in[73] & in[199]); 
    assign layer_0[17] = ~(in[117] ^ in[130]); 
    assign layer_0[18] = ~in[147] | (in[106] & in[147]); 
    assign layer_0[19] = in[203] & ~in[66]; 
    assign layer_0[20] = ~(in[110] ^ in[108]); 
    assign layer_0[21] = ~in[120] | (in[204] & in[120]); 
    assign layer_0[22] = ~(in[200] ^ in[196]); 
    assign layer_0[23] = ~in[57] | (in[57] & in[198]); 
    assign layer_0[24] = ~in[109]; 
    assign layer_0[25] = ~(in[70] | in[165]); 
    assign layer_0[26] = ~(in[87] | in[99]); 
    assign layer_0[27] = ~(in[214] | in[76]); 
    assign layer_0[28] = in[101] | in[197]; 
    assign layer_0[29] = in[230] & ~in[21]; 
    assign layer_0[30] = ~(in[143] | in[5]); 
    assign layer_0[31] = ~(in[198] ^ in[200]); 
    assign layer_0[32] = in[217] & ~in[39]; 
    assign layer_0[33] = in[22] | in[84]; 
    assign layer_0[34] = ~in[186] | (in[186] & in[105]); 
    assign layer_0[35] = in[29] | in[235]; 
    assign layer_0[36] = ~(in[20] ^ in[7]); 
    assign layer_0[37] = in[89] | in[105]; 
    assign layer_0[38] = in[55] ^ in[106]; 
    assign layer_0[39] = ~(in[37] ^ in[68]); 
    assign layer_0[40] = ~(in[31] | in[130]); 
    assign layer_0[41] = in[136]; 
    assign layer_0[42] = in[42]; 
    assign layer_0[43] = in[158] & ~in[103]; 
    assign layer_0[44] = ~(in[183] ^ in[121]); 
    assign layer_0[45] = in[234]; 
    assign layer_0[46] = ~(in[182] ^ in[164]); 
    assign layer_0[47] = ~(in[63] ^ in[95]); 
    assign layer_0[48] = in[180] ^ in[182]; 
    assign layer_0[49] = in[171] | in[59]; 
    assign layer_0[50] = in[152]; 
    assign layer_0[51] = in[145] ^ in[196]; 
    assign layer_0[52] = ~(in[158] | in[62]); 
    assign layer_0[53] = in[121] & ~in[147]; 
    assign layer_0[54] = in[134] & ~in[140]; 
    assign layer_0[55] = ~(in[76] ^ in[45]); 
    assign layer_0[56] = in[145] | in[159]; 
    assign layer_0[57] = ~(in[182] ^ in[146]); 
    assign layer_0[58] = in[92] ^ in[148]; 
    assign layer_0[59] = ~in[138] | (in[138] & in[152]); 
    assign layer_0[60] = ~(in[123] | in[99]); 
    assign layer_0[61] = ~(in[29] ^ in[63]); 
    assign layer_0[62] = ~(in[194] ^ in[218]); 
    assign layer_0[63] = in[90] ^ in[9]; 
    assign layer_0[64] = in[136] & ~in[37]; 
    assign layer_0[65] = ~(in[135] ^ in[164]); 
    assign layer_0[66] = in[142]; 
    assign layer_0[67] = ~(in[76] & in[29]); 
    assign layer_0[68] = ~(in[83] | in[113]); 
    assign layer_0[69] = in[130] ^ in[41]; 
    assign layer_0[70] = ~(in[159] ^ in[230]); 
    assign layer_0[71] = in[122] ^ in[154]; 
    assign layer_0[72] = in[207] ^ in[30]; 
    assign layer_0[73] = ~(in[84] ^ in[70]); 
    assign layer_0[74] = ~in[101] | (in[40] & in[101]); 
    assign layer_0[75] = in[182] ^ in[230]; 
    assign layer_0[76] = in[46] ^ in[94]; 
    assign layer_0[77] = ~(in[103] ^ in[134]); 
    assign layer_0[78] = ~(in[230] ^ in[215]); 
    assign layer_0[79] = in[141] ^ in[154]; 
    assign layer_0[80] = in[103] | in[123]; 
    assign layer_0[81] = ~in[100] | (in[150] & in[100]); 
    assign layer_0[82] = in[241] ^ in[46]; 
    assign layer_0[83] = in[199] & in[234]; 
    assign layer_0[84] = ~(in[118] ^ in[148]); 
    assign layer_0[85] = ~in[90] | (in[70] & in[90]); 
    assign layer_0[86] = ~(in[4] | in[193]); 
    assign layer_0[87] = ~(in[117] ^ in[140]); 
    assign layer_0[88] = ~in[95]; 
    assign layer_0[89] = ~(in[37] ^ in[89]); 
    assign layer_0[90] = ~(in[245] | in[55]); 
    assign layer_0[91] = in[83] | in[52]; 
    assign layer_0[92] = in[181] ^ in[105]; 
    assign layer_0[93] = in[95] ^ in[62]; 
    assign layer_0[94] = in[181] ^ in[164]; 
    assign layer_0[95] = ~(in[119] | in[151]); 
    assign layer_0[96] = ~(in[175] ^ in[194]); 
    assign layer_0[97] = ~(in[79] ^ in[221]); 
    assign layer_0[98] = in[118] | in[103]; 
    assign layer_0[99] = in[58] & ~in[92]; 
    assign layer_0[100] = ~(in[93] ^ in[167]); 
    assign layer_0[101] = ~(in[95] ^ in[58]); 
    assign layer_0[102] = ~(in[126] | in[109]); 
    assign layer_0[103] = ~in[212]; 
    assign layer_0[104] = in[220] | in[142]; 
    assign layer_0[105] = in[11] | in[207]; 
    assign layer_0[106] = ~(in[212] ^ in[198]); 
    assign layer_0[107] = in[171] | in[202]; 
    assign layer_0[108] = in[214] ^ in[167]; 
    assign layer_0[109] = ~in[66] | (in[119] & in[66]); 
    assign layer_0[110] = ~(in[28] | in[220]); 
    assign layer_0[111] = in[199] ^ in[133]; 
    assign layer_0[112] = ~in[27]; 
    assign layer_0[113] = in[92]; 
    assign layer_0[114] = ~in[151]; 
    assign layer_0[115] = in[217]; 
    assign layer_0[116] = ~(in[53] | in[22]); 
    assign layer_0[117] = in[150] | in[165]; 
    assign layer_0[118] = in[173] | in[13]; 
    assign layer_0[119] = in[108] | in[165]; 
    assign layer_0[120] = in[182] & ~in[6]; 
    assign layer_0[121] = in[153] ^ in[217]; 
    assign layer_0[122] = in[86]; 
    assign layer_0[123] = in[218] & ~in[171]; 
    assign layer_0[124] = ~in[74] | (in[74] & in[194]); 
    assign layer_0[125] = in[183] | in[148]; 
    assign layer_0[126] = in[148] | in[51]; 
    assign layer_0[127] = ~(in[118] ^ in[52]); 
    assign layer_0[128] = ~(in[132] | in[37]); 
    assign layer_0[129] = ~in[57] | (in[93] & in[57]); 
    assign layer_0[130] = ~(in[29] ^ in[46]); 
    assign layer_0[131] = ~(in[236] | in[142]); 
    assign layer_0[132] = in[206] ^ in[175]; 
    assign layer_0[133] = ~(in[71] ^ in[36]); 
    assign layer_0[134] = in[137]; 
    assign layer_0[135] = ~(in[35] | in[193]); 
    assign layer_0[136] = ~in[54]; 
    assign layer_0[137] = in[198] | in[198]; 
    assign layer_0[138] = in[137] & ~in[47]; 
    assign layer_0[139] = ~(in[79] ^ in[104]); 
    assign layer_0[140] = in[138] & ~in[157]; 
    assign layer_0[141] = ~(in[179] | in[43]); 
    assign layer_0[142] = in[235] ^ in[59]; 
    assign layer_0[143] = in[200] | in[28]; 
    assign layer_0[144] = in[137] & ~in[156]; 
    assign layer_0[145] = ~(in[210] | in[27]); 
    assign layer_0[146] = ~(in[130] ^ in[116]); 
    assign layer_0[147] = ~(in[105] ^ in[140]); 
    assign layer_0[148] = ~(in[101] ^ in[99]); 
    assign layer_0[149] = in[10] ^ in[30]; 
    assign layer_0[150] = ~in[125]; 
    assign layer_0[151] = in[162] ^ in[153]; 
    assign layer_0[152] = in[90]; 
    assign layer_0[153] = ~in[203] | (in[203] & in[80]); 
    assign layer_0[154] = in[40] & ~in[198]; 
    assign layer_0[155] = in[114] | in[89]; 
    assign layer_0[156] = ~(in[174] | in[173]); 
    assign layer_0[157] = ~in[180] | (in[178] & in[180]); 
    assign layer_0[158] = ~in[163]; 
    assign layer_0[159] = ~(in[185] | in[86]); 
    assign layer_0[160] = ~in[122]; 
    assign layer_0[161] = ~in[182] | (in[182] & in[78]); 
    assign layer_0[162] = ~in[61]; 
    assign layer_0[163] = ~in[105] | (in[105] & in[152]); 
    assign layer_0[164] = ~(in[55] | in[218]); 
    assign layer_0[165] = in[59] & ~in[248]; 
    assign layer_0[166] = in[198] ^ in[151]; 
    assign layer_0[167] = in[199] & ~in[132]; 
    assign layer_0[168] = ~(in[29] | in[184]); 
    assign layer_0[169] = ~in[244]; 
    assign layer_0[170] = in[88]; 
    assign layer_0[171] = in[167]; 
    assign layer_0[172] = in[119] ^ in[150]; 
    assign layer_0[173] = in[21] ^ in[25]; 
    assign layer_0[174] = in[131] ^ in[137]; 
    assign layer_0[175] = ~(in[77] | in[44]); 
    assign layer_0[176] = ~(in[7] | in[6]); 
    assign layer_0[177] = in[152] & ~in[219]; 
    assign layer_0[178] = in[149] ^ in[180]; 
    assign layer_0[179] = ~(in[90] ^ in[123]); 
    assign layer_0[180] = ~(in[213] | in[116]); 
    assign layer_0[181] = in[252] | in[152]; 
    assign layer_0[182] = ~in[137]; 
    assign layer_0[183] = ~in[90] | (in[90] & in[136]); 
    assign layer_0[184] = in[116] | in[210]; 
    assign layer_0[185] = in[105]; 
    assign layer_0[186] = ~(in[202] | in[233]); 
    assign layer_0[187] = ~(in[61] | in[245]); 
    assign layer_0[188] = ~(in[99] | in[94]); 
    assign layer_0[189] = ~(in[151] ^ in[211]); 
    assign layer_0[190] = in[29] | in[61]; 
    assign layer_0[191] = in[218] & ~in[81]; 
    assign layer_0[192] = in[179] ^ in[199]; 
    assign layer_0[193] = in[170]; 
    assign layer_0[194] = ~(in[21] | in[152]); 
    assign layer_0[195] = ~in[99] | (in[99] & in[105]); 
    assign layer_0[196] = ~(in[54] | in[235]); 
    assign layer_0[197] = in[237] | in[169]; 
    assign layer_0[198] = in[168] & ~in[117]; 
    assign layer_0[199] = ~(in[213] ^ in[159]); 
    assign layer_0[200] = ~(in[79] ^ in[243]); 
    assign layer_0[201] = ~(in[146] ^ in[163]); 
    assign layer_0[202] = in[187] | in[92]; 
    assign layer_0[203] = in[131] ^ in[133]; 
    assign layer_0[204] = ~(in[78] ^ in[98]); 
    assign layer_0[205] = in[165] ^ in[185]; 
    assign layer_0[206] = in[151] & ~in[245]; 
    assign layer_0[207] = ~in[148] | (in[148] & in[59]); 
    assign layer_0[208] = in[154] ^ in[59]; 
    assign layer_0[209] = ~(in[120] ^ in[151]); 
    assign layer_0[210] = ~(in[88] | in[117]); 
    assign layer_0[211] = ~(in[136] | in[137]); 
    assign layer_0[212] = in[84] ^ in[181]; 
    assign layer_0[213] = ~(in[204] | in[212]); 
    assign layer_0[214] = ~in[133]; 
    assign layer_0[215] = ~(in[236] ^ in[21]); 
    assign layer_0[216] = ~(in[138] | in[105]); 
    assign layer_0[217] = in[127] ^ in[141]; 
    assign layer_0[218] = ~in[247]; 
    assign layer_0[219] = ~(in[75] | in[133]); 
    assign layer_0[220] = ~in[123]; 
    assign layer_0[221] = in[235]; 
    assign layer_0[222] = in[126] & ~in[138]; 
    assign layer_0[223] = in[56] ^ in[103]; 
    assign layer_0[224] = in[72] ^ in[86]; 
    assign layer_0[225] = ~(in[83] ^ in[104]); 
    assign layer_0[226] = in[164] ^ in[40]; 
    assign layer_0[227] = ~in[134] | (in[172] & in[134]); 
    assign layer_0[228] = in[193] ^ in[36]; 
    assign layer_0[229] = ~(in[199] ^ in[43]); 
    assign layer_0[230] = ~in[243]; 
    assign layer_0[231] = ~(in[247] | in[231]); 
    assign layer_0[232] = in[207] ^ in[159]; 
    assign layer_0[233] = in[120] | in[111]; 
    assign layer_0[234] = ~(in[222] ^ in[65]); 
    assign layer_0[235] = in[130] | in[103]; 
    assign layer_0[236] = in[103] ^ in[56]; 
    assign layer_0[237] = in[25] ^ in[28]; 
    assign layer_0[238] = in[232] | in[143]; 
    assign layer_0[239] = in[192] | in[36]; 
    assign layer_0[240] = in[122] | in[157]; 
    assign layer_0[241] = ~(in[178] ^ in[180]); 
    assign layer_0[242] = in[132]; 
    assign layer_0[243] = ~(in[71] | in[89]); 
    assign layer_0[244] = in[131]; 
    assign layer_0[245] = ~(in[194] ^ in[119]); 
    assign layer_0[246] = ~(in[56] ^ in[95]); 
    assign layer_0[247] = ~in[154] | (in[154] & in[118]); 
    assign layer_0[248] = in[90] & in[140]; 
    assign layer_0[249] = ~(in[36] ^ in[68]); 
    assign layer_0[250] = in[214] & ~in[30]; 
    assign layer_0[251] = in[102] ^ in[87]; 
    assign layer_0[252] = in[210]; 
    assign layer_0[253] = in[171]; 
    assign layer_0[254] = ~(in[143] | in[131]); 
    assign layer_0[255] = in[139] & in[138]; 
    assign layer_0[256] = ~in[227]; 
    assign layer_0[257] = in[149] ^ in[152]; 
    assign layer_0[258] = in[115] & ~in[117]; 
    assign layer_0[259] = ~in[89]; 
    assign layer_0[260] = in[153] & ~in[203]; 
    assign layer_0[261] = ~(in[237] ^ in[248]); 
    assign layer_0[262] = ~in[74]; 
    assign layer_0[263] = ~(in[155] ^ in[182]); 
    assign layer_0[264] = in[203] ^ in[180]; 
    assign layer_0[265] = ~(in[107] ^ in[75]); 
    assign layer_0[266] = ~(in[119] ^ in[150]); 
    assign layer_0[267] = in[184] ^ in[138]; 
    assign layer_0[268] = ~(in[121] | in[155]); 
    assign layer_0[269] = in[57] | in[42]; 
    assign layer_0[270] = ~in[181]; 
    assign layer_0[271] = ~(in[153] ^ in[35]); 
    assign layer_0[272] = ~in[232]; 
    assign layer_0[273] = in[59] & ~in[116]; 
    assign layer_0[274] = ~(in[103] | in[117]); 
    assign layer_0[275] = in[235]; 
    assign layer_0[276] = ~in[46] | (in[46] & in[56]); 
    assign layer_0[277] = ~(in[133] | in[164]); 
    assign layer_0[278] = ~in[213] | (in[213] & in[227]); 
    assign layer_0[279] = in[231] ^ in[241]; 
    assign layer_0[280] = in[46] | in[138]; 
    assign layer_0[281] = in[87] ^ in[90]; 
    assign layer_0[282] = ~(in[124] ^ in[163]); 
    assign layer_0[283] = in[78] | in[43]; 
    assign layer_0[284] = ~(in[213] | in[55]); 
    assign layer_0[285] = in[111] | in[158]; 
    assign layer_0[286] = ~in[248]; 
    assign layer_0[287] = in[213] ^ in[177]; 
    assign layer_0[288] = ~(in[73] | in[75]); 
    assign layer_0[289] = in[147] & ~in[76]; 
    assign layer_0[290] = ~(in[173] ^ in[89]); 
    assign layer_0[291] = ~in[155]; 
    assign layer_0[292] = in[221] | in[175]; 
    assign layer_0[293] = ~(in[220] | in[131]); 
    assign layer_0[294] = in[177] ^ in[8]; 
    assign layer_0[295] = in[105] & ~in[101]; 
    assign layer_0[296] = ~in[216] | (in[247] & in[216]); 
    assign layer_0[297] = in[70] | in[185]; 
    assign layer_0[298] = ~in[185] | (in[185] & in[213]); 
    assign layer_0[299] = ~(in[39] | in[55]); 
    assign layer_0[300] = 1'b1; 
    assign layer_0[301] = ~in[136]; 
    assign layer_0[302] = in[98] ^ in[245]; 
    assign layer_0[303] = in[170] ^ in[103]; 
    assign layer_0[304] = in[154]; 
    assign layer_0[305] = ~in[163] | (in[163] & in[54]); 
    assign layer_0[306] = in[164] ^ in[166]; 
    assign layer_0[307] = in[241] & ~in[232]; 
    assign layer_0[308] = in[174] | in[35]; 
    assign layer_0[309] = ~(in[83] ^ in[58]); 
    assign layer_0[310] = in[162] ^ in[62]; 
    assign layer_0[311] = ~(in[22] ^ in[24]); 
    assign layer_0[312] = ~(in[19] ^ in[7]); 
    assign layer_0[313] = ~in[137] | (in[90] & in[137]); 
    assign layer_0[314] = in[35]; 
    assign layer_0[315] = in[114] ^ in[37]; 
    assign layer_0[316] = ~(in[124] | in[122]); 
    assign layer_0[317] = in[8] ^ in[177]; 
    assign layer_0[318] = in[29] & ~in[170]; 
    assign layer_0[319] = ~in[133] | (in[68] & in[133]); 
    assign layer_0[320] = ~in[221]; 
    assign layer_0[321] = ~(in[109] ^ in[111]); 
    assign layer_0[322] = ~in[130] | (in[130] & in[120]); 
    assign layer_0[323] = in[198] & ~in[100]; 
    assign layer_0[324] = in[109] | in[211]; 
    assign layer_0[325] = ~(in[21] | in[163]); 
    assign layer_0[326] = in[114] ^ in[41]; 
    assign layer_0[327] = in[93] ^ in[46]; 
    assign layer_0[328] = in[79] & ~in[123]; 
    assign layer_0[329] = in[134] ^ in[102]; 
    assign layer_0[330] = ~in[104] | (in[156] & in[104]); 
    assign layer_0[331] = in[91] & ~in[216]; 
    assign layer_0[332] = ~(in[87] ^ in[228]); 
    assign layer_0[333] = in[118] ^ in[172]; 
    assign layer_0[334] = ~in[136] | (in[136] & in[116]); 
    assign layer_0[335] = in[232] ^ in[184]; 
    assign layer_0[336] = ~in[58]; 
    assign layer_0[337] = ~(in[163] | in[233]); 
    assign layer_0[338] = in[187] | in[50]; 
    assign layer_0[339] = in[182] & ~in[42]; 
    assign layer_0[340] = in[234]; 
    assign layer_0[341] = ~(in[206] | in[126]); 
    assign layer_0[342] = in[123] | in[178]; 
    assign layer_0[343] = ~in[169] | (in[169] & in[211]); 
    assign layer_0[344] = ~(in[146] | in[133]); 
    assign layer_0[345] = ~(in[113] | in[125]); 
    assign layer_0[346] = ~in[40]; 
    assign layer_0[347] = ~in[52] | (in[42] & in[52]); 
    assign layer_0[348] = ~in[137]; 
    assign layer_0[349] = in[27]; 
    assign layer_0[350] = ~(in[78] | in[139]); 
    assign layer_0[351] = ~in[182] | (in[244] & in[182]); 
    assign layer_0[352] = in[231] | in[54]; 
    assign layer_0[353] = in[241]; 
    assign layer_0[354] = in[67] ^ in[185]; 
    assign layer_0[355] = in[54] ^ in[7]; 
    assign layer_0[356] = ~(in[143] | in[199]); 
    assign layer_0[357] = in[230] & ~in[244]; 
    assign layer_0[358] = ~(in[43] & in[126]); 
    assign layer_0[359] = in[178] ^ in[137]; 
    assign layer_0[360] = ~in[150] | (in[157] & in[150]); 
    assign layer_0[361] = ~in[86] | (in[151] & in[86]); 
    assign layer_0[362] = in[77] ^ in[73]; 
    assign layer_0[363] = in[99]; 
    assign layer_0[364] = in[62] ^ in[44]; 
    assign layer_0[365] = in[104] | in[183]; 
    assign layer_0[366] = in[138] ^ in[121]; 
    assign layer_0[367] = in[52] ^ in[82]; 
    assign layer_0[368] = in[245] ^ in[214]; 
    assign layer_0[369] = in[78] | in[86]; 
    assign layer_0[370] = ~(in[127] ^ in[117]); 
    assign layer_0[371] = in[187] ^ in[235]; 
    assign layer_0[372] = ~(in[102] & in[251]); 
    assign layer_0[373] = in[233]; 
    assign layer_0[374] = in[76] | in[124]; 
    assign layer_0[375] = in[120] & ~in[101]; 
    assign layer_0[376] = ~in[149] | (in[149] & in[212]); 
    assign layer_0[377] = ~(in[93] & in[109]); 
    assign layer_0[378] = ~(in[146] | in[78]); 
    assign layer_0[379] = ~in[169] | (in[169] & in[234]); 
    assign layer_0[380] = in[66] ^ in[105]; 
    assign layer_0[381] = in[198] ^ in[229]; 
    assign layer_0[382] = in[187] ^ in[55]; 
    assign layer_0[383] = ~(in[229] | in[214]); 
    assign layer_0[384] = in[196] ^ in[182]; 
    assign layer_0[385] = in[117] & ~in[197]; 
    assign layer_0[386] = in[143] | in[116]; 
    assign layer_0[387] = ~(in[166] ^ in[197]); 
    assign layer_0[388] = ~(in[100] ^ in[105]); 
    assign layer_0[389] = in[194] | in[135]; 
    assign layer_0[390] = in[143] | in[158]; 
    assign layer_0[391] = in[93] ^ in[111]; 
    assign layer_0[392] = ~in[70] | (in[103] & in[70]); 
    assign layer_0[393] = in[93] ^ in[56]; 
    assign layer_0[394] = in[244] ^ in[95]; 
    assign layer_0[395] = ~(in[98] ^ in[84]); 
    assign layer_0[396] = ~(in[53] ^ in[66]); 
    assign layer_0[397] = in[88] & in[89]; 
    assign layer_0[398] = in[152] | in[161]; 
    assign layer_0[399] = in[192] | in[204]; 
    assign layer_0[400] = in[179] & ~in[137]; 
    assign layer_0[401] = ~(in[117] ^ in[102]); 
    assign layer_0[402] = ~in[251] | (in[188] & in[251]); 
    assign layer_0[403] = ~in[101] | (in[101] & in[83]); 
    assign layer_0[404] = in[52] | in[155]; 
    assign layer_0[405] = in[100] | in[191]; 
    assign layer_0[406] = in[214] | in[159]; 
    assign layer_0[407] = ~(in[70] ^ in[38]); 
    assign layer_0[408] = ~(in[8] | in[21]); 
    assign layer_0[409] = ~(in[213] & in[211]); 
    assign layer_0[410] = ~(in[45] | in[59]); 
    assign layer_0[411] = in[165] ^ in[148]; 
    assign layer_0[412] = in[115] | in[98]; 
    assign layer_0[413] = ~in[168]; 
    assign layer_0[414] = ~(in[172] | in[198]); 
    assign layer_0[415] = ~(in[75] ^ in[24]); 
    assign layer_0[416] = in[91] ^ in[51]; 
    assign layer_0[417] = ~in[163]; 
    assign layer_0[418] = in[154] ^ in[186]; 
    assign layer_0[419] = in[228] | in[120]; 
    assign layer_0[420] = ~in[36]; 
    assign layer_0[421] = ~(in[196] ^ in[131]); 
    assign layer_0[422] = in[92] | in[247]; 
    assign layer_0[423] = in[182] | in[164]; 
    assign layer_0[424] = ~in[137]; 
    assign layer_0[425] = in[72] ^ in[24]; 
    assign layer_0[426] = in[251] | in[67]; 
    assign layer_0[427] = in[149] & ~in[245]; 
    assign layer_0[428] = ~in[217] | (in[217] & in[249]); 
    assign layer_0[429] = ~(in[169] ^ in[216]); 
    assign layer_0[430] = in[186] & ~in[117]; 
    assign layer_0[431] = in[75]; 
    assign layer_0[432] = in[121] & ~in[167]; 
    assign layer_0[433] = in[115] | in[183]; 
    assign layer_0[434] = in[109] | in[106]; 
    assign layer_0[435] = in[168] & ~in[92]; 
    assign layer_0[436] = in[115] | in[172]; 
    assign layer_0[437] = in[147] ^ in[165]; 
    assign layer_0[438] = in[251] ^ in[220]; 
    assign layer_0[439] = in[216] ^ in[249]; 
    assign layer_0[440] = in[46] | in[30]; 
    assign layer_0[441] = ~in[166] | (in[166] & in[43]); 
    assign layer_0[442] = ~(in[78] ^ in[80]); 
    assign layer_0[443] = in[168] | in[170]; 
    assign layer_0[444] = ~(in[152] | in[136]); 
    assign layer_0[445] = ~(in[26] ^ in[52]); 
    assign layer_0[446] = in[41] | in[117]; 
    assign layer_0[447] = ~(in[77] ^ in[7]); 
    assign layer_0[448] = ~(in[97] | in[99]); 
    assign layer_0[449] = ~(in[47] | in[145]); 
    assign layer_0[450] = ~in[55] | (in[168] & in[55]); 
    assign layer_0[451] = ~(in[135] ^ in[152]); 
    assign layer_0[452] = in[45] ^ in[79]; 
    assign layer_0[453] = ~in[117] | (in[8] & in[117]); 
    assign layer_0[454] = in[184] ^ in[152]; 
    assign layer_0[455] = in[103] | in[168]; 
    assign layer_0[456] = in[183] & ~in[85]; 
    assign layer_0[457] = ~(in[102] ^ in[97]); 
    assign layer_0[458] = in[111] ^ in[49]; 
    assign layer_0[459] = in[108] ^ in[90]; 
    assign layer_0[460] = ~(in[72] ^ in[76]); 
    assign layer_0[461] = ~(in[36] | in[152]); 
    assign layer_0[462] = ~(in[101] ^ in[98]); 
    assign layer_0[463] = ~in[75]; 
    assign layer_0[464] = ~in[90]; 
    assign layer_0[465] = ~in[87]; 
    assign layer_0[466] = in[27] | in[95]; 
    assign layer_0[467] = ~in[137]; 
    assign layer_0[468] = in[179] | in[58]; 
    assign layer_0[469] = in[87] ^ in[114]; 
    assign layer_0[470] = ~in[230] | (in[183] & in[230]); 
    assign layer_0[471] = ~(in[43] ^ in[108]); 
    assign layer_0[472] = ~in[121] | (in[187] & in[121]); 
    assign layer_0[473] = ~(in[191] | in[207]); 
    assign layer_0[474] = in[57] & ~in[8]; 
    assign layer_0[475] = ~(in[219] | in[164]); 
    assign layer_0[476] = ~in[70] | (in[70] & in[101]); 
    assign layer_0[477] = in[216]; 
    assign layer_0[478] = ~in[108] | (in[108] & in[178]); 
    assign layer_0[479] = ~in[119] | (in[167] & in[119]); 
    assign layer_0[480] = in[166] ^ in[69]; 
    assign layer_0[481] = in[231] ^ in[135]; 
    assign layer_0[482] = in[26] & ~in[150]; 
    assign layer_0[483] = in[180] | in[198]; 
    assign layer_0[484] = ~(in[40] | in[114]); 
    assign layer_0[485] = ~in[152] | (in[152] & in[99]); 
    assign layer_0[486] = ~in[195]; 
    assign layer_0[487] = in[9] & ~in[109]; 
    assign layer_0[488] = in[88] | in[210]; 
    assign layer_0[489] = in[133] & in[95]; 
    assign layer_0[490] = ~in[181] | (in[181] & in[53]); 
    assign layer_0[491] = ~(in[103] ^ in[71]); 
    assign layer_0[492] = ~in[145]; 
    assign layer_0[493] = in[104] ^ in[74]; 
    assign layer_0[494] = in[78] | in[151]; 
    assign layer_0[495] = in[51] ^ in[197]; 
    assign layer_0[496] = in[130] | in[244]; 
    assign layer_0[497] = ~in[107] | (in[107] & in[94]); 
    assign layer_0[498] = in[118] & ~in[162]; 
    assign layer_0[499] = ~(in[145] | in[159]); 
    assign layer_0[500] = ~(in[87] ^ in[179]); 
    assign layer_0[501] = in[165] & ~in[78]; 
    assign layer_0[502] = in[101] | in[100]; 
    assign layer_0[503] = in[106] ^ in[23]; 
    assign layer_0[504] = ~(in[166] ^ in[198]); 
    assign layer_0[505] = in[23] ^ in[69]; 
    assign layer_0[506] = ~in[156] | (in[156] & in[194]); 
    assign layer_0[507] = ~(in[241] ^ in[223]); 
    assign layer_0[508] = ~(in[61] | in[74]); 
    assign layer_0[509] = ~(in[85] | in[106]); 
    assign layer_0[510] = ~(in[21] | in[195]); 
    assign layer_0[511] = in[181] ^ in[124]; 
    assign layer_0[512] = ~(in[198] ^ in[196]); 
    assign layer_0[513] = in[58] ^ in[29]; 
    assign layer_0[514] = in[90] ^ in[108]; 
    assign layer_0[515] = ~(in[210] | in[54]); 
    assign layer_0[516] = in[155] | in[52]; 
    assign layer_0[517] = ~(in[218] ^ in[140]); 
    assign layer_0[518] = ~(in[107] ^ in[46]); 
    assign layer_0[519] = ~in[155] | (in[155] & in[213]); 
    assign layer_0[520] = in[57]; 
    assign layer_0[521] = in[58] & ~in[62]; 
    assign layer_0[522] = ~(in[163] | in[156]); 
    assign layer_0[523] = ~in[156]; 
    assign layer_0[524] = ~(in[122] ^ in[137]); 
    assign layer_0[525] = ~in[53]; 
    assign layer_0[526] = in[43] ^ in[76]; 
    assign layer_0[527] = in[150] ^ in[148]; 
    assign layer_0[528] = in[201] ^ in[70]; 
    assign layer_0[529] = ~(in[29] & in[76]); 
    assign layer_0[530] = ~(in[63] | in[188]); 
    assign layer_0[531] = in[170] ^ in[102]; 
    assign layer_0[532] = in[85] & ~in[71]; 
    assign layer_0[533] = in[230] | in[41]; 
    assign layer_0[534] = in[188] | in[190]; 
    assign layer_0[535] = ~in[232] | (in[201] & in[232]); 
    assign layer_0[536] = in[218] & ~in[109]; 
    assign layer_0[537] = ~(in[119] | in[135]); 
    assign layer_0[538] = ~in[121] | (in[127] & in[121]); 
    assign layer_0[539] = ~in[118] | (in[91] & in[118]); 
    assign layer_0[540] = in[163]; 
    assign layer_0[541] = ~(in[50] | in[129]); 
    assign layer_0[542] = in[245]; 
    assign layer_0[543] = ~in[152] | (in[213] & in[152]); 
    assign layer_0[544] = ~in[63]; 
    assign layer_0[545] = ~(in[165] ^ in[245]); 
    assign layer_0[546] = in[181] ^ in[183]; 
    assign layer_0[547] = ~in[148]; 
    assign layer_0[548] = in[183] ^ in[139]; 
    assign layer_0[549] = ~(in[250] | in[169]); 
    assign layer_0[550] = ~(in[50] ^ in[208]); 
    assign layer_0[551] = ~in[183] | (in[183] & in[27]); 
    assign layer_0[552] = ~(in[171] ^ in[121]); 
    assign layer_0[553] = in[232] ^ in[195]; 
    assign layer_0[554] = in[87]; 
    assign layer_0[555] = ~in[134] | (in[136] & in[134]); 
    assign layer_0[556] = ~in[134]; 
    assign layer_0[557] = ~(in[69] ^ in[188]); 
    assign layer_0[558] = in[92] ^ in[116]; 
    assign layer_0[559] = in[71] ^ in[103]; 
    assign layer_0[560] = in[218] & ~in[237]; 
    assign layer_0[561] = ~(in[228] ^ in[51]); 
    assign layer_0[562] = in[158] ^ in[196]; 
    assign layer_0[563] = in[117] ^ in[146]; 
    assign layer_0[564] = in[147]; 
    assign layer_0[565] = in[86] ^ in[100]; 
    assign layer_0[566] = ~(in[182] & in[196]); 
    assign layer_0[567] = in[171] | in[138]; 
    assign layer_0[568] = in[131] | in[130]; 
    assign layer_0[569] = in[22] ^ in[36]; 
    assign layer_0[570] = ~in[137] | (in[137] & in[53]); 
    assign layer_0[571] = ~(in[193] | in[218]); 
    assign layer_0[572] = in[87] & ~in[206]; 
    assign layer_0[573] = 1'b1; 
    assign layer_0[574] = ~(in[172] ^ in[170]); 
    assign layer_0[575] = ~in[135] | (in[135] & in[55]); 
    assign layer_0[576] = in[156] | in[241]; 
    assign layer_0[577] = in[139] ^ in[134]; 
    assign layer_0[578] = in[115] ^ in[132]; 
    assign layer_0[579] = in[133] | in[132]; 
    assign layer_0[580] = in[41] & ~in[155]; 
    assign layer_0[581] = in[202]; 
    assign layer_0[582] = ~in[29]; 
    assign layer_0[583] = ~in[42] | (in[42] & in[167]); 
    assign layer_0[584] = ~(in[88] ^ in[41]); 
    assign layer_0[585] = in[225] | in[152]; 
    assign layer_0[586] = in[116] ^ in[102]; 
    assign layer_0[587] = in[219]; 
    assign layer_0[588] = ~(in[141] ^ in[82]); 
    assign layer_0[589] = in[114] ^ in[100]; 
    assign layer_0[590] = ~in[12]; 
    assign layer_0[591] = ~(in[85] | in[100]); 
    assign layer_0[592] = ~(in[210] ^ in[245]); 
    assign layer_0[593] = in[95]; 
    assign layer_0[594] = ~(in[84] ^ in[87]); 
    assign layer_0[595] = in[197] ^ in[178]; 
    assign layer_0[596] = in[146] & ~in[103]; 
    assign layer_0[597] = ~(in[85] | in[214]); 
    assign layer_0[598] = ~(in[169] ^ in[130]); 
    assign layer_0[599] = ~(in[147] | in[118]); 
    assign layer_0[600] = ~(in[59] ^ in[90]); 
    assign layer_0[601] = ~(in[40] ^ in[9]); 
    assign layer_0[602] = in[171] ^ in[124]; 
    assign layer_0[603] = in[104]; 
    assign layer_0[604] = ~(in[182] ^ in[151]); 
    assign layer_0[605] = ~(in[201] ^ in[232]); 
    assign layer_0[606] = in[131] & ~in[197]; 
    assign layer_0[607] = ~in[137] | (in[203] & in[137]); 
    assign layer_0[608] = ~(in[197] | in[196]); 
    assign layer_0[609] = ~(in[241] ^ in[11]); 
    assign layer_0[610] = in[243] ^ in[196]; 
    assign layer_0[611] = in[87] ^ in[104]; 
    assign layer_0[612] = in[72] & ~in[59]; 
    assign layer_0[613] = in[142] | in[24]; 
    assign layer_0[614] = ~(in[174] | in[228]); 
    assign layer_0[615] = in[113] | in[114]; 
    assign layer_0[616] = ~(in[90] ^ in[23]); 
    assign layer_0[617] = in[140]; 
    assign layer_0[618] = ~in[186]; 
    assign layer_0[619] = ~in[9]; 
    assign layer_0[620] = ~in[186]; 
    assign layer_0[621] = in[119] | in[137]; 
    assign layer_0[622] = in[199] & ~in[186]; 
    assign layer_0[623] = in[147] & ~in[43]; 
    assign layer_0[624] = in[124]; 
    assign layer_0[625] = in[185] ^ in[167]; 
    assign layer_0[626] = in[123] & in[136]; 
    assign layer_0[627] = ~in[213] | (in[213] & in[87]); 
    assign layer_0[628] = ~in[70] | (in[164] & in[70]); 
    assign layer_0[629] = in[153]; 
    assign layer_0[630] = ~(in[164] ^ in[134]); 
    assign layer_0[631] = ~(in[23] ^ in[58]); 
    assign layer_0[632] = ~(in[195] | in[145]); 
    assign layer_0[633] = ~in[212] | (in[212] & in[51]); 
    assign layer_0[634] = in[213] & ~in[46]; 
    assign layer_0[635] = ~(in[85] ^ in[243]); 
    assign layer_0[636] = in[159] | in[8]; 
    assign layer_0[637] = ~(in[78] ^ in[31]); 
    assign layer_0[638] = ~in[219]; 
    assign layer_0[639] = in[29] | in[4]; 
    assign layer_0[640] = in[94] | in[132]; 
    assign layer_0[641] = in[226] ^ in[100]; 
    assign layer_0[642] = ~in[209]; 
    assign layer_0[643] = ~(in[178] ^ in[213]); 
    assign layer_0[644] = in[168] & ~in[126]; 
    assign layer_0[645] = ~(in[141] | in[140]); 
    assign layer_0[646] = ~(in[164] | in[183]); 
    assign layer_0[647] = in[236] ^ in[111]; 
    assign layer_0[648] = ~in[105] | (in[179] & in[105]); 
    assign layer_0[649] = ~(in[184] | in[227]); 
    assign layer_0[650] = ~(in[247] ^ in[79]); 
    assign layer_0[651] = in[56] | in[140]; 
    assign layer_0[652] = ~in[196]; 
    assign layer_0[653] = ~(in[171] | in[154]); 
    assign layer_0[654] = ~in[8] | (in[54] & in[8]); 
    assign layer_0[655] = in[210]; 
    assign layer_0[656] = ~in[61] | (in[61] & in[103]); 
    assign layer_0[657] = ~(in[107] ^ in[183]); 
    assign layer_0[658] = ~(in[34] | in[176]); 
    assign layer_0[659] = ~(in[66] ^ in[35]); 
    assign layer_0[660] = in[165] ^ in[163]; 
    assign layer_0[661] = ~in[156]; 
    assign layer_0[662] = ~in[92]; 
    assign layer_0[663] = ~(in[11] ^ in[83]); 
    assign layer_0[664] = ~in[227]; 
    assign layer_0[665] = in[29] | in[146]; 
    assign layer_0[666] = ~in[106]; 
    assign layer_0[667] = ~(in[94] ^ in[77]); 
    assign layer_0[668] = ~(in[98] | in[162]); 
    assign layer_0[669] = ~in[151]; 
    assign layer_0[670] = in[109] & ~in[47]; 
    assign layer_0[671] = ~in[199] | (in[245] & in[199]); 
    assign layer_0[672] = in[119] | in[214]; 
    assign layer_0[673] = ~(in[102] ^ in[116]); 
    assign layer_0[674] = in[71] & ~in[42]; 
    assign layer_0[675] = ~in[171]; 
    assign layer_0[676] = in[131]; 
    assign layer_0[677] = ~(in[211] | in[251]); 
    assign layer_0[678] = ~in[82]; 
    assign layer_0[679] = ~in[159] | (in[134] & in[159]); 
    assign layer_0[680] = in[132] | in[76]; 
    assign layer_0[681] = ~(in[71] ^ in[24]); 
    assign layer_0[682] = in[109] | in[126]; 
    assign layer_0[683] = in[242] | in[174]; 
    assign layer_0[684] = ~(in[82] ^ in[68]); 
    assign layer_0[685] = in[86] & ~in[143]; 
    assign layer_0[686] = ~in[172] | (in[172] & in[186]); 
    assign layer_0[687] = in[212] & ~in[166]; 
    assign layer_0[688] = ~(in[210] ^ in[57]); 
    assign layer_0[689] = in[106] ^ in[88]; 
    assign layer_0[690] = in[210] ^ in[6]; 
    assign layer_0[691] = ~(in[126] ^ in[134]); 
    assign layer_0[692] = ~(in[140] & in[80]); 
    assign layer_0[693] = in[57] ^ in[104]; 
    assign layer_0[694] = in[118] ^ in[116]; 
    assign layer_0[695] = in[27] | in[10]; 
    assign layer_0[696] = ~(in[75] ^ in[73]); 
    assign layer_0[697] = in[98] ^ in[83]; 
    assign layer_0[698] = in[212] & ~in[121]; 
    assign layer_0[699] = in[106] & ~in[133]; 
    assign layer_0[700] = ~(in[162] | in[164]); 
    assign layer_0[701] = in[136] & ~in[115]; 
    assign layer_0[702] = in[181] & ~in[106]; 
    assign layer_0[703] = in[57] ^ in[55]; 
    assign layer_0[704] = ~in[138] | (in[184] & in[138]); 
    assign layer_0[705] = in[238] | in[113]; 
    assign layer_0[706] = ~(in[53] ^ in[5]); 
    assign layer_0[707] = ~in[140]; 
    assign layer_0[708] = ~(in[130] | in[242]); 
    assign layer_0[709] = in[194] ^ in[165]; 
    assign layer_0[710] = in[117] & ~in[34]; 
    assign layer_0[711] = in[212] | in[62]; 
    assign layer_0[712] = ~(in[40] ^ in[72]); 
    assign layer_0[713] = ~(in[34] ^ in[65]); 
    assign layer_0[714] = in[228] | in[213]; 
    assign layer_0[715] = in[103] ^ in[189]; 
    assign layer_0[716] = ~(in[68] ^ in[86]); 
    assign layer_0[717] = in[49] | in[5]; 
    assign layer_0[718] = in[191] | in[243]; 
    assign layer_0[719] = ~in[120] | (in[120] & in[124]); 
    assign layer_0[720] = in[10] | in[86]; 
    assign layer_0[721] = ~(in[27] | in[232]); 
    assign layer_0[722] = in[163] | in[74]; 
    assign layer_0[723] = ~(in[44] ^ in[42]); 
    assign layer_0[724] = in[157] ^ in[234]; 
    assign layer_0[725] = ~in[245]; 
    assign layer_0[726] = in[11]; 
    assign layer_0[727] = in[55] ^ in[56]; 
    assign layer_0[728] = ~(in[172] ^ in[101]); 
    assign layer_0[729] = ~(in[143] | in[194]); 
    assign layer_0[730] = ~(in[233] ^ in[202]); 
    assign layer_0[731] = in[168]; 
    assign layer_0[732] = ~(in[149] ^ in[146]); 
    assign layer_0[733] = ~(in[147] ^ in[134]); 
    assign layer_0[734] = in[174] & in[174]; 
    assign layer_0[735] = in[118] & ~in[99]; 
    assign layer_0[736] = in[187]; 
    assign layer_0[737] = ~in[136] | (in[155] & in[136]); 
    assign layer_0[738] = ~(in[183] ^ in[89]); 
    assign layer_0[739] = ~in[42] | (in[42] & in[131]); 
    assign layer_0[740] = in[165] & ~in[167]; 
    assign layer_0[741] = ~(in[186] ^ in[234]); 
    assign layer_0[742] = in[166] ^ in[149]; 
    assign layer_0[743] = ~(in[183] | in[180]); 
    assign layer_0[744] = ~in[217] | (in[157] & in[217]); 
    assign layer_0[745] = ~(in[131] | in[168]); 
    assign layer_0[746] = in[165] ^ in[202]; 
    assign layer_0[747] = ~(in[87] ^ in[55]); 
    assign layer_0[748] = in[170] ^ in[37]; 
    assign layer_0[749] = in[90] ^ in[108]; 
    assign layer_0[750] = in[150] & ~in[25]; 
    assign layer_0[751] = ~in[78]; 
    assign layer_0[752] = ~(in[99] | in[163]); 
    assign layer_0[753] = in[101] ^ in[115]; 
    assign layer_0[754] = in[164] ^ in[182]; 
    assign layer_0[755] = ~(in[75] ^ in[77]); 
    assign layer_0[756] = ~in[187] | (in[187] & in[137]); 
    assign layer_0[757] = ~(in[167] | in[7]); 
    assign layer_0[758] = ~in[38] | (in[38] & in[7]); 
    assign layer_0[759] = ~(in[54] ^ in[103]); 
    assign layer_0[760] = in[68] & ~in[137]; 
    assign layer_0[761] = ~in[170]; 
    assign layer_0[762] = in[150] & ~in[105]; 
    assign layer_0[763] = in[156]; 
    assign layer_0[764] = in[8] & ~in[165]; 
    assign layer_0[765] = ~in[126]; 
    assign layer_0[766] = in[249] ^ in[87]; 
    assign layer_0[767] = in[74]; 
    assign layer_0[768] = ~in[182] | (in[216] & in[182]); 
    assign layer_0[769] = in[23] ^ in[121]; 
    assign layer_0[770] = ~(in[251] | in[151]); 
    assign layer_0[771] = in[209] ^ in[156]; 
    assign layer_0[772] = ~(in[44] ^ in[194]); 
    assign layer_0[773] = ~(in[102] ^ in[70]); 
    assign layer_0[774] = ~in[130]; 
    assign layer_0[775] = in[147] | in[103]; 
    assign layer_0[776] = ~(in[203] | in[172]); 
    assign layer_0[777] = ~in[138] | (in[138] & in[143]); 
    assign layer_0[778] = in[152] & ~in[117]; 
    assign layer_0[779] = in[189] ^ in[141]; 
    assign layer_0[780] = in[244] | in[204]; 
    assign layer_0[781] = in[120] ^ in[4]; 
    assign layer_0[782] = in[182] ^ in[184]; 
    assign layer_0[783] = in[41] ^ in[156]; 
    assign layer_0[784] = ~in[230] | (in[61] & in[230]); 
    assign layer_0[785] = in[137] & ~in[234]; 
    assign layer_0[786] = in[220] & ~in[117]; 
    assign layer_0[787] = in[154] ^ in[36]; 
    assign layer_0[788] = ~(in[228] ^ in[182]); 
    assign layer_0[789] = in[85]; 
    assign layer_0[790] = in[188] | in[194]; 
    assign layer_0[791] = in[214] & ~in[107]; 
    assign layer_0[792] = ~(in[184] | in[137]); 
    assign layer_0[793] = ~(in[6] ^ in[228]); 
    assign layer_0[794] = ~(in[135] | in[5]); 
    assign layer_0[795] = in[245] ^ in[198]; 
    assign layer_0[796] = in[170] ^ in[183]; 
    assign layer_0[797] = in[67] & ~in[54]; 
    assign layer_0[798] = ~(in[149] | in[90]); 
    assign layer_0[799] = ~in[183] | (in[183] & in[210]); 
    assign layer_0[800] = ~(in[91] ^ in[77]); 
    assign layer_0[801] = in[141]; 
    assign layer_0[802] = ~in[180]; 
    assign layer_0[803] = in[84] | in[72]; 
    assign layer_0[804] = ~(in[140] | in[203]); 
    assign layer_0[805] = in[89] ^ in[211]; 
    assign layer_0[806] = ~(in[183] ^ in[230]); 
    assign layer_0[807] = ~(in[36] ^ in[22]); 
    assign layer_0[808] = in[120] | in[113]; 
    assign layer_0[809] = ~(in[191] ^ in[62]); 
    assign layer_0[810] = in[99] ^ in[117]; 
    assign layer_0[811] = ~(in[96] | in[66]); 
    assign layer_0[812] = in[197]; 
    assign layer_0[813] = in[136] ^ in[199]; 
    assign layer_0[814] = ~in[162] | (in[162] & in[122]); 
    assign layer_0[815] = in[134] ^ in[119]; 
    assign layer_0[816] = ~(in[228] ^ in[168]); 
    assign layer_0[817] = ~(in[116] & in[220]); 
    assign layer_0[818] = ~(in[149] | in[116]); 
    assign layer_0[819] = ~(in[104] | in[95]); 
    assign layer_0[820] = ~(in[156] ^ in[58]); 
    assign layer_0[821] = in[164]; 
    assign layer_0[822] = ~(in[69] | in[51]); 
    assign layer_0[823] = ~(in[243] ^ in[223]); 
    assign layer_0[824] = ~(in[211] ^ in[246]); 
    assign layer_0[825] = in[188] ^ in[219]; 
    assign layer_0[826] = in[59] ^ in[122]; 
    assign layer_0[827] = in[90]; 
    assign layer_0[828] = in[140] ^ in[242]; 
    assign layer_0[829] = ~in[72] | (in[157] & in[72]); 
    assign layer_0[830] = in[54] ^ in[85]; 
    assign layer_0[831] = in[23] | in[102]; 
    assign layer_0[832] = in[71] | in[182]; 
    assign layer_0[833] = in[73] | in[172]; 
    assign layer_0[834] = in[171]; 
    assign layer_0[835] = ~in[85]; 
    assign layer_0[836] = in[23] & ~in[53]; 
    assign layer_0[837] = ~(in[190] | in[184]); 
    assign layer_0[838] = in[23] ^ in[71]; 
    assign layer_0[839] = in[217] ^ in[135]; 
    assign layer_0[840] = in[214] & ~in[210]; 
    assign layer_0[841] = in[134] & ~in[181]; 
    assign layer_0[842] = ~in[93]; 
    assign layer_0[843] = ~in[95]; 
    assign layer_0[844] = in[119] & ~in[221]; 
    assign layer_0[845] = ~in[104]; 
    assign layer_0[846] = in[50] | in[249]; 
    assign layer_0[847] = in[234] | in[193]; 
    assign layer_0[848] = in[92] ^ in[55]; 
    assign layer_0[849] = ~(in[250] | in[217]); 
    assign layer_0[850] = ~(in[102] | in[63]); 
    assign layer_0[851] = in[47] ^ in[209]; 
    assign layer_0[852] = in[108] & ~in[158]; 
    assign layer_0[853] = ~(in[111] | in[5]); 
    assign layer_0[854] = ~in[232] | (in[211] & in[232]); 
    assign layer_0[855] = ~(in[5] | in[34]); 
    assign layer_0[856] = in[135] ^ in[96]; 
    assign layer_0[857] = in[202] & ~in[141]; 
    assign layer_0[858] = in[95] ^ in[8]; 
    assign layer_0[859] = in[41]; 
    assign layer_0[860] = in[136]; 
    assign layer_0[861] = in[183]; 
    assign layer_0[862] = ~(in[110] ^ in[108]); 
    assign layer_0[863] = in[235] ^ in[186]; 
    assign layer_0[864] = ~(in[24] ^ in[70]); 
    assign layer_0[865] = ~in[29] | (in[29] & in[229]); 
    assign layer_0[866] = ~in[28]; 
    assign layer_0[867] = in[54] & ~in[251]; 
    assign layer_0[868] = in[85] ^ in[68]; 
    assign layer_0[869] = ~(in[163] ^ in[162]); 
    assign layer_0[870] = ~in[199] | (in[42] & in[199]); 
    assign layer_0[871] = ~(in[109] ^ in[83]); 
    assign layer_0[872] = ~in[47]; 
    assign layer_0[873] = ~in[34]; 
    assign layer_0[874] = in[183] ^ in[124]; 
    assign layer_0[875] = in[170] & ~in[205]; 
    assign layer_0[876] = in[118]; 
    assign layer_0[877] = in[110] | in[98]; 
    assign layer_0[878] = in[113] | in[41]; 
    assign layer_0[879] = ~(in[92] | in[26]); 
    assign layer_0[880] = in[170]; 
    assign layer_0[881] = in[246] | in[212]; 
    assign layer_0[882] = ~(in[95] | in[75]); 
    assign layer_0[883] = ~(in[115] ^ in[175]); 
    assign layer_0[884] = in[220] | in[236]; 
    assign layer_0[885] = ~(in[127] ^ in[175]); 
    assign layer_0[886] = in[41] & ~in[39]; 
    assign layer_0[887] = in[186] & ~in[54]; 
    assign layer_0[888] = in[146] | in[148]; 
    assign layer_0[889] = ~(in[230] ^ in[198]); 
    assign layer_0[890] = in[77] & in[245]; 
    assign layer_0[891] = ~(in[89] ^ in[99]); 
    assign layer_0[892] = ~(in[93] | in[41]); 
    assign layer_0[893] = ~(in[221] ^ in[79]); 
    assign layer_0[894] = ~(in[134] | in[196]); 
    assign layer_0[895] = in[114] | in[174]; 
    assign layer_0[896] = in[117]; 
    assign layer_0[897] = in[70] & ~in[57]; 
    assign layer_0[898] = in[102] ^ in[99]; 
    assign layer_0[899] = ~(in[196] ^ in[218]); 
    assign layer_0[900] = ~(in[91] | in[78]); 
    assign layer_0[901] = in[95] | in[47]; 
    assign layer_0[902] = in[181]; 
    assign layer_0[903] = ~(in[236] ^ in[250]); 
    assign layer_0[904] = ~in[85] | (in[60] & in[85]); 
    assign layer_0[905] = in[213] & ~in[50]; 
    assign layer_0[906] = in[163]; 
    assign layer_0[907] = in[237] ^ in[205]; 
    assign layer_0[908] = ~(in[90] ^ in[146]); 
    assign layer_0[909] = in[137]; 
    assign layer_0[910] = in[90]; 
    assign layer_0[911] = ~(in[8] ^ in[177]); 
    assign layer_0[912] = ~(in[236] ^ in[151]); 
    assign layer_0[913] = in[181]; 
    assign layer_0[914] = ~(in[103] | in[120]); 
    assign layer_0[915] = in[152] | in[148]; 
    assign layer_0[916] = in[182] | in[165]; 
    assign layer_0[917] = ~(in[57] ^ in[26]); 
    assign layer_0[918] = in[104] ^ in[147]; 
    assign layer_0[919] = in[90] ^ in[108]; 
    assign layer_0[920] = ~(in[87] ^ in[40]); 
    assign layer_0[921] = ~(in[249] ^ in[59]); 
    assign layer_0[922] = ~in[102] | (in[102] & in[180]); 
    assign layer_0[923] = in[184] & in[131]; 
    assign layer_0[924] = in[149] ^ in[147]; 
    assign layer_0[925] = ~(in[39] ^ in[71]); 
    assign layer_0[926] = in[114] ^ in[79]; 
    assign layer_0[927] = in[83] ^ in[12]; 
    assign layer_0[928] = ~(in[102] | in[89]); 
    assign layer_0[929] = in[230] & ~in[10]; 
    assign layer_0[930] = ~(in[105] ^ in[137]); 
    assign layer_0[931] = ~(in[247] | in[241]); 
    assign layer_0[932] = in[228] ^ in[198]; 
    assign layer_0[933] = ~(in[112] | in[165]); 
    assign layer_0[934] = ~(in[78] ^ in[148]); 
    assign layer_0[935] = in[214] | in[228]; 
    assign layer_0[936] = in[141]; 
    assign layer_0[937] = ~in[138] | (in[138] & in[196]); 
    assign layer_0[938] = in[167] & ~in[107]; 
    assign layer_0[939] = ~in[94] | (in[94] & in[157]); 
    assign layer_0[940] = in[50] | in[202]; 
    assign layer_0[941] = ~(in[202] ^ in[234]); 
    assign layer_0[942] = in[116] & ~in[24]; 
    assign layer_0[943] = in[201] ^ in[143]; 
    assign layer_0[944] = in[91] & ~in[251]; 
    assign layer_0[945] = ~(in[107] | in[212]); 
    assign layer_0[946] = in[87] ^ in[57]; 
    assign layer_0[947] = in[121] & ~in[157]; 
    assign layer_0[948] = ~in[88] | (in[38] & in[88]); 
    assign layer_0[949] = in[166] | in[167]; 
    assign layer_0[950] = in[158] ^ in[217]; 
    assign layer_0[951] = ~(in[116] | in[102]); 
    assign layer_0[952] = ~(in[207] | in[186]); 
    assign layer_0[953] = in[37] ^ in[83]; 
    assign layer_0[954] = in[44] | in[136]; 
    assign layer_0[955] = ~in[39] | (in[62] & in[39]); 
    assign layer_0[956] = in[249] ^ in[233]; 
    assign layer_0[957] = in[221]; 
    assign layer_0[958] = ~(in[21] | in[193]); 
    assign layer_0[959] = in[13] | in[30]; 
    assign layer_0[960] = ~in[108] | (in[158] & in[108]); 
    assign layer_0[961] = in[73] ^ in[43]; 
    assign layer_0[962] = ~(in[205] | in[195]); 
    assign layer_0[963] = in[183] ^ in[120]; 
    assign layer_0[964] = ~(in[177] | in[83]); 
    assign layer_0[965] = in[60] ^ in[94]; 
    assign layer_0[966] = ~in[201] | (in[74] & in[201]); 
    assign layer_0[967] = ~(in[198] | in[188]); 
    assign layer_0[968] = ~(in[116] | in[147]); 
    assign layer_0[969] = in[198] | in[197]; 
    assign layer_0[970] = in[46] ^ in[108]; 
    assign layer_0[971] = in[53] & ~in[189]; 
    assign layer_0[972] = ~in[118]; 
    assign layer_0[973] = in[101] | in[211]; 
    assign layer_0[974] = in[132] ^ in[134]; 
    assign layer_0[975] = in[15]; 
    assign layer_0[976] = ~(in[38] ^ in[195]); 
    assign layer_0[977] = in[216] | in[22]; 
    assign layer_0[978] = in[149] & ~in[55]; 
    assign layer_0[979] = ~(in[88] ^ in[91]); 
    assign layer_0[980] = in[123] ^ in[91]; 
    assign layer_0[981] = in[174] | in[137]; 
    assign layer_0[982] = ~in[187] | (in[134] & in[187]); 
    assign layer_0[983] = in[221] ^ in[13]; 
    assign layer_0[984] = in[78]; 
    assign layer_0[985] = in[196] | in[54]; 
    assign layer_0[986] = ~in[230] | (in[218] & in[230]); 
    assign layer_0[987] = ~(in[94] ^ in[65]); 
    assign layer_0[988] = ~(in[75] | in[133]); 
    assign layer_0[989] = ~in[181] | (in[243] & in[181]); 
    assign layer_0[990] = ~(in[205] ^ in[138]); 
    assign layer_0[991] = in[117] ^ in[171]; 
    assign layer_0[992] = in[91] ^ in[60]; 
    assign layer_0[993] = ~(in[21] | in[192]); 
    assign layer_0[994] = ~(in[146] ^ in[62]); 
    assign layer_0[995] = in[181]; 
    assign layer_0[996] = in[245]; 
    assign layer_0[997] = ~(in[94] ^ in[76]); 
    assign layer_0[998] = in[69] & in[72]; 
    assign layer_0[999] = ~(in[189] ^ in[220]); 
    assign layer_0[1000] = ~(in[8] & in[43]); 
    assign layer_0[1001] = ~(in[151] | in[117]); 
    assign layer_0[1002] = ~in[149] | (in[105] & in[149]); 
    assign layer_0[1003] = ~in[98]; 
    assign layer_0[1004] = in[172] | in[36]; 
    assign layer_0[1005] = in[107]; 
    assign layer_0[1006] = in[187] & in[168]; 
    assign layer_0[1007] = in[92] ^ in[45]; 
    assign layer_0[1008] = ~(in[166] ^ in[164]); 
    assign layer_0[1009] = ~in[169]; 
    assign layer_0[1010] = in[158] ^ in[205]; 
    assign layer_0[1011] = in[54] | in[38]; 
    assign layer_0[1012] = ~(in[187] ^ in[38]); 
    assign layer_0[1013] = in[117] & in[173]; 
    assign layer_0[1014] = ~(in[41] ^ in[71]); 
    assign layer_0[1015] = ~in[217] | (in[217] & in[211]); 
    assign layer_0[1016] = in[70] ^ in[84]; 
    assign layer_0[1017] = ~in[131]; 
    assign layer_0[1018] = ~(in[197] | in[50]); 
    assign layer_0[1019] = in[249] & ~in[246]; 
    assign layer_0[1020] = ~(in[242] | in[157]); 
    assign layer_0[1021] = ~(in[109] ^ in[69]); 
    assign layer_0[1022] = in[140] | in[72]; 
    assign layer_0[1023] = in[151] ^ in[69]; 
    assign layer_0[1024] = in[173] ^ in[205]; 
    assign layer_0[1025] = in[60] | in[65]; 
    assign layer_0[1026] = ~(in[212] ^ in[93]); 
    assign layer_0[1027] = in[216]; 
    assign layer_0[1028] = in[78] | in[134]; 
    assign layer_0[1029] = in[131] ^ in[170]; 
    assign layer_0[1030] = ~(in[148] ^ in[146]); 
    assign layer_0[1031] = in[120]; 
    assign layer_0[1032] = in[251] | in[74]; 
    assign layer_0[1033] = in[235]; 
    assign layer_0[1034] = in[148] ^ in[130]; 
    assign layer_0[1035] = ~(in[108] | in[25]); 
    assign layer_0[1036] = in[211] ^ in[151]; 
    assign layer_0[1037] = ~(in[84] | in[194]); 
    assign layer_0[1038] = ~(in[82] ^ in[117]); 
    assign layer_0[1039] = in[101] & ~in[73]; 
    assign layer_0[1040] = in[20] | in[233]; 
    assign layer_0[1041] = ~(in[246] | in[79]); 
    assign layer_0[1042] = in[166]; 
    assign layer_0[1043] = in[102] ^ in[91]; 
    assign layer_0[1044] = in[28] & ~in[106]; 
    assign layer_0[1045] = in[55] ^ in[185]; 
    assign layer_0[1046] = ~in[229]; 
    assign layer_0[1047] = ~in[37] | (in[199] & in[37]); 
    assign layer_0[1048] = in[78] ^ in[77]; 
    assign layer_0[1049] = in[8] & ~in[235]; 
    assign layer_0[1050] = in[131]; 
    assign layer_0[1051] = ~(in[219] ^ in[173]); 
    assign layer_0[1052] = in[166] | in[167]; 
    assign layer_0[1053] = in[167] & ~in[86]; 
    assign layer_0[1054] = in[156] & ~in[120]; 
    assign layer_0[1055] = ~in[123] | (in[184] & in[123]); 
    assign layer_0[1056] = ~(in[130] ^ in[226]); 
    assign layer_0[1057] = in[90] | in[92]; 
    assign layer_0[1058] = in[84]; 
    assign layer_0[1059] = ~(in[124] ^ in[107]); 
    assign layer_0[1060] = in[227] | in[205]; 
    assign layer_0[1061] = in[93] ^ in[216]; 
    assign layer_0[1062] = in[126] | in[12]; 
    assign layer_0[1063] = in[198] | in[212]; 
    assign layer_0[1064] = in[75] & ~in[235]; 
    assign layer_0[1065] = ~(in[82] ^ in[135]); 
    assign layer_0[1066] = in[166] | in[164]; 
    assign layer_0[1067] = in[56] ^ in[85]; 
    assign layer_0[1068] = ~in[188] | (in[188] & in[183]); 
    assign layer_0[1069] = ~(in[166] ^ in[50]); 
    assign layer_0[1070] = in[62] ^ in[221]; 
    assign layer_0[1071] = in[24] & ~in[150]; 
    assign layer_0[1072] = ~in[104] | (in[104] & in[141]); 
    assign layer_0[1073] = ~(in[9] | in[63]); 
    assign layer_0[1074] = ~in[23] | (in[110] & in[23]); 
    assign layer_0[1075] = ~(in[132] ^ in[119]); 
    assign layer_0[1076] = ~(in[19] | in[151]); 
    assign layer_0[1077] = ~in[200]; 
    assign layer_0[1078] = in[69] | in[243]; 
    assign layer_0[1079] = in[154] & ~in[27]; 
    assign layer_0[1080] = ~in[93] | (in[93] & in[117]); 
    assign layer_0[1081] = in[143] | in[21]; 
    assign layer_0[1082] = in[172] | in[89]; 
    assign layer_0[1083] = ~(in[91] ^ in[93]); 
    assign layer_0[1084] = ~(in[244] ^ in[96]); 
    assign layer_0[1085] = in[181] & ~in[178]; 
    assign layer_0[1086] = in[24] ^ in[56]; 
    assign layer_0[1087] = ~(in[101] | in[100]); 
    assign layer_0[1088] = in[228] & ~in[88]; 
    assign layer_0[1089] = ~(in[237] | in[11]); 
    assign layer_0[1090] = in[150]; 
    assign layer_0[1091] = in[194] & ~in[111]; 
    assign layer_0[1092] = in[135]; 
    assign layer_0[1093] = in[209] ^ in[11]; 
    assign layer_0[1094] = in[28] | in[41]; 
    assign layer_0[1095] = in[153] ^ in[119]; 
    assign layer_0[1096] = ~in[207]; 
    assign layer_0[1097] = ~in[52] | (in[74] & in[52]); 
    assign layer_0[1098] = in[102] & ~in[84]; 
    assign layer_0[1099] = ~in[30]; 
    assign layer_0[1100] = in[103] ^ in[36]; 
    assign layer_0[1101] = ~in[123] | (in[58] & in[123]); 
    assign layer_0[1102] = ~(in[197] ^ in[83]); 
    assign layer_0[1103] = in[138] & ~in[68]; 
    assign layer_0[1104] = ~(in[115] ^ in[102]); 
    assign layer_0[1105] = in[123] | in[155]; 
    assign layer_0[1106] = ~in[200] | (in[100] & in[200]); 
    assign layer_0[1107] = ~in[59] | (in[203] & in[59]); 
    assign layer_0[1108] = in[154] ^ in[119]; 
    assign layer_0[1109] = ~in[165] | (in[165] & in[62]); 
    assign layer_0[1110] = ~(in[215] | in[248]); 
    assign layer_0[1111] = in[138] ^ in[187]; 
    assign layer_0[1112] = in[66] ^ in[172]; 
    assign layer_0[1113] = in[9] & ~in[42]; 
    assign layer_0[1114] = ~(in[205] | in[21]); 
    assign layer_0[1115] = in[35] & in[221]; 
    assign layer_0[1116] = ~in[214] | (in[214] & in[107]); 
    assign layer_0[1117] = ~(in[199] ^ in[214]); 
    assign layer_0[1118] = in[79] ^ in[46]; 
    assign layer_0[1119] = in[94] ^ in[39]; 
    assign layer_0[1120] = ~(in[186] ^ in[199]); 
    assign layer_0[1121] = in[132] & ~in[218]; 
    assign layer_0[1122] = in[91] & ~in[119]; 
    assign layer_0[1123] = ~(in[25] | in[106]); 
    assign layer_0[1124] = ~(in[105] ^ in[153]); 
    assign layer_0[1125] = in[103] & ~in[75]; 
    assign layer_0[1126] = ~in[88]; 
    assign layer_0[1127] = in[107] & in[105]; 
    assign layer_0[1128] = ~in[24]; 
    assign layer_0[1129] = ~(in[126] | in[124]); 
    assign layer_0[1130] = in[230]; 
    assign layer_0[1131] = in[126] & ~in[136]; 
    assign layer_0[1132] = in[206] ^ in[195]; 
    assign layer_0[1133] = in[148] | in[147]; 
    assign layer_0[1134] = ~(in[227] | in[199]); 
    assign layer_0[1135] = ~in[39] | (in[39] & in[170]); 
    assign layer_0[1136] = ~in[71] | (in[155] & in[71]); 
    assign layer_0[1137] = ~in[24] | (in[60] & in[24]); 
    assign layer_0[1138] = in[21] | in[226]; 
    assign layer_0[1139] = ~(in[93] ^ in[91]); 
    assign layer_0[1140] = ~(in[55] & in[115]); 
    assign layer_0[1141] = in[226] ^ in[131]; 
    assign layer_0[1142] = in[133] ^ in[28]; 
    assign layer_0[1143] = ~in[109]; 
    assign layer_0[1144] = ~(in[249] ^ in[236]); 
    assign layer_0[1145] = in[151] & in[101]; 
    assign layer_0[1146] = ~(in[21] | in[59]); 
    assign layer_0[1147] = in[12] ^ in[83]; 
    assign layer_0[1148] = ~in[100] | (in[211] & in[100]); 
    assign layer_0[1149] = in[72] & ~in[123]; 
    assign layer_0[1150] = ~(in[92] | in[107]); 
    assign layer_0[1151] = in[27] & ~in[122]; 
    assign layer_0[1152] = in[71] ^ in[90]; 
    assign layer_0[1153] = in[200] ^ in[218]; 
    assign layer_0[1154] = in[82] ^ in[95]; 
    assign layer_0[1155] = in[114] ^ in[63]; 
    assign layer_0[1156] = in[38] ^ in[203]; 
    assign layer_0[1157] = ~(in[247] | in[249]); 
    assign layer_0[1158] = in[135] ^ in[104]; 
    assign layer_0[1159] = in[11] | in[9]; 
    assign layer_0[1160] = in[88] | in[120]; 
    assign layer_0[1161] = ~(in[204] | in[181]); 
    assign layer_0[1162] = in[71] & ~in[187]; 
    assign layer_0[1163] = ~(in[90] ^ in[201]); 
    assign layer_0[1164] = ~(in[115] ^ in[102]); 
    assign layer_0[1165] = in[196] ^ in[82]; 
    assign layer_0[1166] = in[103]; 
    assign layer_0[1167] = ~(in[235] ^ in[196]); 
    assign layer_0[1168] = in[118] & ~in[123]; 
    assign layer_0[1169] = ~(in[175] | in[162]); 
    assign layer_0[1170] = in[196]; 
    assign layer_0[1171] = in[85] | in[54]; 
    assign layer_0[1172] = ~in[245] | (in[197] & in[245]); 
    assign layer_0[1173] = ~(in[88] | in[177]); 
    assign layer_0[1174] = ~in[24] | (in[74] & in[24]); 
    assign layer_0[1175] = ~(in[105] ^ in[125]); 
    assign layer_0[1176] = in[137] ^ in[105]; 
    assign layer_0[1177] = ~in[181] | (in[23] & in[181]); 
    assign layer_0[1178] = in[197] | in[24]; 
    assign layer_0[1179] = in[76]; 
    assign layer_0[1180] = in[11] & ~in[84]; 
    assign layer_0[1181] = in[70] & ~in[153]; 
    assign layer_0[1182] = ~(in[198] ^ in[169]); 
    assign layer_0[1183] = ~in[153] | (in[153] & in[82]); 
    assign layer_0[1184] = ~(in[142] ^ in[155]); 
    assign layer_0[1185] = ~(in[135] ^ in[43]); 
    assign layer_0[1186] = ~in[88] | (in[42] & in[88]); 
    assign layer_0[1187] = in[196] & ~in[220]; 
    assign layer_0[1188] = in[90] ^ in[108]; 
    assign layer_0[1189] = in[98] ^ in[99]; 
    assign layer_0[1190] = in[27] & ~in[56]; 
    assign layer_0[1191] = ~(in[168] | in[150]); 
    assign layer_0[1192] = ~(in[151] | in[126]); 
    assign layer_0[1193] = ~in[227]; 
    assign layer_0[1194] = in[51] & ~in[55]; 
    assign layer_0[1195] = ~(in[155] | in[177]); 
    assign layer_0[1196] = ~(in[227] | in[88]); 
    assign layer_0[1197] = ~in[166] | (in[243] & in[166]); 
    assign layer_0[1198] = in[177] ^ in[209]; 
    assign layer_0[1199] = ~(in[110] ^ in[92]); 
    assign layer_0[1200] = ~(in[46] ^ in[107]); 
    assign layer_0[1201] = ~(in[204] | in[247]); 
    assign layer_0[1202] = in[123] & ~in[142]; 
    assign layer_0[1203] = ~(in[36] ^ in[22]); 
    assign layer_0[1204] = ~in[126] | (in[112] & in[126]); 
    assign layer_0[1205] = in[46] ^ in[215]; 
    assign layer_0[1206] = ~(in[85] ^ in[188]); 
    assign layer_0[1207] = in[59] ^ in[91]; 
    assign layer_0[1208] = in[71] ^ in[25]; 
    assign layer_0[1209] = in[171] | in[154]; 
    assign layer_0[1210] = ~in[70]; 
    assign layer_0[1211] = ~in[27] | (in[27] & in[84]); 
    assign layer_0[1212] = in[109] ^ in[123]; 
    assign layer_0[1213] = in[124]; 
    assign layer_0[1214] = ~in[129]; 
    assign layer_0[1215] = ~in[147]; 
    assign layer_0[1216] = ~(in[170] | in[163]); 
    assign layer_0[1217] = ~(in[235] | in[94]); 
    assign layer_0[1218] = ~(in[11] ^ in[161]); 
    assign layer_0[1219] = ~(in[190] | in[205]); 
    assign layer_0[1220] = ~(in[94] ^ in[106]); 
    assign layer_0[1221] = in[56] ^ in[24]; 
    assign layer_0[1222] = ~(in[181] | in[236]); 
    assign layer_0[1223] = ~(in[74] ^ in[211]); 
    assign layer_0[1224] = ~(in[118] ^ in[88]); 
    assign layer_0[1225] = ~(in[47] | in[193]); 
    assign layer_0[1226] = ~in[152] | (in[109] & in[152]); 
    assign layer_0[1227] = ~in[182] | (in[182] & in[247]); 
    assign layer_0[1228] = in[116] & ~in[37]; 
    assign layer_0[1229] = ~(in[54] ^ in[105]); 
    assign layer_0[1230] = in[152] ^ in[105]; 
    assign layer_0[1231] = ~(in[200] | in[90]); 
    assign layer_0[1232] = ~(in[106] ^ in[141]); 
    assign layer_0[1233] = in[61] ^ in[44]; 
    assign layer_0[1234] = ~(in[78] ^ in[45]); 
    assign layer_0[1235] = ~(in[150] | in[126]); 
    assign layer_0[1236] = ~(in[183] | in[21]); 
    assign layer_0[1237] = ~(in[232] ^ in[183]); 
    assign layer_0[1238] = ~(in[94] | in[173]); 
    assign layer_0[1239] = in[92] & ~in[151]; 
    assign layer_0[1240] = in[41] ^ in[72]; 
    assign layer_0[1241] = ~(in[170] & in[236]); 
    assign layer_0[1242] = ~in[235] | (in[235] & in[248]); 
    assign layer_0[1243] = ~(in[198] ^ in[228]); 
    assign layer_0[1244] = in[189] | in[210]; 
    assign layer_0[1245] = in[170] ^ in[54]; 
    assign layer_0[1246] = in[114] | in[98]; 
    assign layer_0[1247] = in[198]; 
    assign layer_0[1248] = ~(in[109] ^ in[82]); 
    assign layer_0[1249] = ~(in[170] ^ in[148]); 
    assign layer_0[1250] = in[122] ^ in[156]; 
    assign layer_0[1251] = in[196] ^ in[220]; 
    assign layer_0[1252] = ~(in[5] | in[143]); 
    assign layer_0[1253] = ~(in[182] ^ in[180]); 
    assign layer_0[1254] = in[77] ^ in[53]; 
    assign layer_0[1255] = in[210] ^ in[247]; 
    assign layer_0[1256] = ~in[154]; 
    assign layer_0[1257] = ~in[209]; 
    assign layer_0[1258] = ~(in[72] & in[131]); 
    assign layer_0[1259] = in[86] & in[190]; 
    assign layer_0[1260] = in[242] ^ in[210]; 
    assign layer_0[1261] = ~(in[42] | in[117]); 
    assign layer_0[1262] = in[250] ^ in[129]; 
    assign layer_0[1263] = in[245]; 
    assign layer_0[1264] = ~(in[72] ^ in[44]); 
    assign layer_0[1265] = ~in[206]; 
    assign layer_0[1266] = ~(in[148] | in[168]); 
    assign layer_0[1267] = ~in[210]; 
    assign layer_0[1268] = in[106]; 
    assign layer_0[1269] = ~(in[156] ^ in[198]); 
    assign layer_0[1270] = in[103] ^ in[113]; 
    assign layer_0[1271] = in[196] | in[236]; 
    assign layer_0[1272] = in[133] & ~in[68]; 
    assign layer_0[1273] = in[183] ^ in[186]; 
    assign layer_0[1274] = ~in[126] | (in[135] & in[126]); 
    assign layer_0[1275] = ~(in[109] | in[93]); 
    assign layer_0[1276] = in[76] ^ in[25]; 
    assign layer_0[1277] = ~in[74] | (in[136] & in[74]); 
    assign layer_0[1278] = in[194] | in[250]; 
    assign layer_0[1279] = in[13] | in[30]; 
    assign layer_0[1280] = ~in[163] | (in[163] & in[194]); 
    assign layer_0[1281] = ~in[136]; 
    assign layer_0[1282] = ~(in[206] ^ in[235]); 
    assign layer_0[1283] = in[193] ^ in[190]; 
    assign layer_0[1284] = ~(in[92] | in[56]); 
    assign layer_0[1285] = in[103]; 
    assign layer_0[1286] = ~in[168] | (in[168] & in[38]); 
    assign layer_0[1287] = in[93]; 
    assign layer_0[1288] = in[178] ^ in[175]; 
    assign layer_0[1289] = ~(in[199] ^ in[148]); 
    assign layer_0[1290] = in[79] ^ in[127]; 
    assign layer_0[1291] = ~(in[103] | in[189]); 
    assign layer_0[1292] = in[194] ^ in[27]; 
    assign layer_0[1293] = in[50] | in[81]; 
    assign layer_0[1294] = in[168]; 
    assign layer_0[1295] = in[71] ^ in[74]; 
    assign layer_0[1296] = in[72]; 
    assign layer_0[1297] = ~(in[147] ^ in[168]); 
    assign layer_0[1298] = ~(in[243] & in[197]); 
    assign layer_0[1299] = ~(in[232] | in[151]); 
    assign layer_0[1300] = in[103] ^ in[58]; 
    assign layer_0[1301] = ~(in[214] | in[94]); 
    assign layer_0[1302] = ~in[119] | (in[119] & in[149]); 
    assign layer_0[1303] = ~(in[60] | in[120]); 
    assign layer_0[1304] = in[237] ^ in[177]; 
    assign layer_0[1305] = in[164] & in[180]; 
    assign layer_0[1306] = in[242] ^ in[185]; 
    assign layer_0[1307] = 1'b0; 
    assign layer_0[1308] = ~(in[152] ^ in[88]); 
    assign layer_0[1309] = ~(in[21] | in[213]); 
    assign layer_0[1310] = in[124] | in[104]; 
    assign layer_0[1311] = ~(in[57] | in[41]); 
    assign layer_0[1312] = ~(in[120] ^ in[98]); 
    assign layer_0[1313] = in[162] ^ in[199]; 
    assign layer_0[1314] = ~(in[172] | in[135]); 
    assign layer_0[1315] = ~(in[179] ^ in[215]); 
    assign layer_0[1316] = ~(in[59] | in[107]); 
    assign layer_0[1317] = ~(in[130] | in[124]); 
    assign layer_0[1318] = ~(in[114] | in[180]); 
    assign layer_0[1319] = in[190] | in[179]; 
    assign layer_0[1320] = ~(in[202] ^ in[251]); 
    assign layer_0[1321] = in[216] | in[232]; 
    assign layer_0[1322] = in[117] | in[163]; 
    assign layer_0[1323] = in[219] | in[219]; 
    assign layer_0[1324] = in[130] & in[115]; 
    assign layer_0[1325] = in[103] & ~in[100]; 
    assign layer_0[1326] = in[149]; 
    assign layer_0[1327] = in[219] ^ in[251]; 
    assign layer_0[1328] = ~(in[148] ^ in[119]); 
    assign layer_0[1329] = in[58]; 
    assign layer_0[1330] = in[206] ^ in[154]; 
    assign layer_0[1331] = ~(in[38] ^ in[41]); 
    assign layer_0[1332] = ~(in[213] ^ in[159]); 
    assign layer_0[1333] = in[220] ^ in[249]; 
    assign layer_0[1334] = ~(in[129] | in[94]); 
    assign layer_0[1335] = ~(in[72] | in[53]); 
    assign layer_0[1336] = ~(in[198] ^ in[244]); 
    assign layer_0[1337] = in[72] ^ in[40]; 
    assign layer_0[1338] = in[137] & ~in[155]; 
    assign layer_0[1339] = in[170]; 
    assign layer_0[1340] = in[214] | in[116]; 
    assign layer_0[1341] = ~(in[186] | in[26]); 
    assign layer_0[1342] = in[89] ^ in[104]; 
    assign layer_0[1343] = in[235] ^ in[209]; 
    assign layer_0[1344] = in[242] & ~in[182]; 
    assign layer_0[1345] = ~(in[95] ^ in[190]); 
    assign layer_0[1346] = in[59] | in[231]; 
    assign layer_0[1347] = ~(in[69] ^ in[52]); 
    assign layer_0[1348] = ~in[90]; 
    assign layer_0[1349] = in[60] | in[200]; 
    assign layer_0[1350] = ~in[126]; 
    assign layer_0[1351] = in[104] ^ in[83]; 
    assign layer_0[1352] = ~(in[37] | in[226]); 
    assign layer_0[1353] = ~(in[155] | in[54]); 
    assign layer_0[1354] = in[171] | in[173]; 
    assign layer_0[1355] = in[34] | in[152]; 
    assign layer_0[1356] = ~(in[235] | in[221]); 
    assign layer_0[1357] = in[198] & ~in[184]; 
    assign layer_0[1358] = ~(in[58] ^ in[90]); 
    assign layer_0[1359] = ~(in[252] ^ in[203]); 
    assign layer_0[1360] = in[179] ^ in[181]; 
    assign layer_0[1361] = in[172] & ~in[87]; 
    assign layer_0[1362] = ~(in[68] | in[151]); 
    assign layer_0[1363] = in[51] ^ in[72]; 
    assign layer_0[1364] = ~in[91]; 
    assign layer_0[1365] = in[38] ^ in[234]; 
    assign layer_0[1366] = ~(in[197] | in[179]); 
    assign layer_0[1367] = ~(in[140] | in[157]); 
    assign layer_0[1368] = ~(in[249] | in[46]); 
    assign layer_0[1369] = in[155] ^ in[52]; 
    assign layer_0[1370] = ~(in[186] & in[155]); 
    assign layer_0[1371] = in[56] ^ in[22]; 
    assign layer_0[1372] = in[150] | in[130]; 
    assign layer_0[1373] = in[89] | in[125]; 
    assign layer_0[1374] = ~(in[118] ^ in[104]); 
    assign layer_0[1375] = in[52] ^ in[186]; 
    assign layer_0[1376] = ~(in[100] ^ in[86]); 
    assign layer_0[1377] = in[74] ^ in[76]; 
    assign layer_0[1378] = in[35] ^ in[137]; 
    assign layer_0[1379] = ~in[214] | (in[120] & in[214]); 
    assign layer_0[1380] = in[91] ^ in[44]; 
    assign layer_0[1381] = in[26] ^ in[75]; 
    assign layer_0[1382] = ~in[40] | (in[149] & in[40]); 
    assign layer_0[1383] = ~(in[164] ^ in[182]); 
    assign layer_0[1384] = ~(in[197] ^ in[195]); 
    assign layer_0[1385] = in[141] ^ in[126]; 
    assign layer_0[1386] = ~in[167] | (in[167] & in[175]); 
    assign layer_0[1387] = ~(in[197] ^ in[143]); 
    assign layer_0[1388] = ~(in[218] ^ in[111]); 
    assign layer_0[1389] = ~(in[170] | in[101]); 
    assign layer_0[1390] = in[169] & ~in[177]; 
    assign layer_0[1391] = ~(in[78] | in[138]); 
    assign layer_0[1392] = ~in[132]; 
    assign layer_0[1393] = ~(in[165] ^ in[250]); 
    assign layer_0[1394] = ~(in[218] | in[101]); 
    assign layer_0[1395] = in[45] | in[20]; 
    assign layer_0[1396] = in[56] | in[79]; 
    assign layer_0[1397] = ~(in[153] & in[170]); 
    assign layer_0[1398] = in[117]; 
    assign layer_0[1399] = in[87] ^ in[220]; 
    assign layer_0[1400] = ~in[131]; 
    assign layer_0[1401] = in[202] & ~in[92]; 
    assign layer_0[1402] = ~in[59] | (in[59] & in[98]); 
    assign layer_0[1403] = ~in[143]; 
    assign layer_0[1404] = in[197] ^ in[228]; 
    assign layer_0[1405] = ~(in[52] ^ in[83]); 
    assign layer_0[1406] = ~in[165] | (in[165] & in[211]); 
    assign layer_0[1407] = ~(in[22] ^ in[70]); 
    assign layer_0[1408] = ~(in[232] | in[196]); 
    assign layer_0[1409] = in[11] | in[207]; 
    assign layer_0[1410] = ~in[147]; 
    assign layer_0[1411] = ~(in[88] ^ in[197]); 
    assign layer_0[1412] = ~in[73]; 
    assign layer_0[1413] = in[167] & ~in[196]; 
    assign layer_0[1414] = ~(in[19] ^ in[208]); 
    assign layer_0[1415] = ~(in[194] ^ in[195]); 
    assign layer_0[1416] = in[70] & ~in[27]; 
    assign layer_0[1417] = ~in[165] | (in[165] & in[107]); 
    assign layer_0[1418] = in[138]; 
    assign layer_0[1419] = in[176] | in[18]; 
    assign layer_0[1420] = ~(in[218] ^ in[187]); 
    assign layer_0[1421] = ~in[151] | (in[218] & in[151]); 
    assign layer_0[1422] = in[167] & in[185]; 
    assign layer_0[1423] = in[181] ^ in[86]; 
    assign layer_0[1424] = in[253]; 
    assign layer_0[1425] = ~(in[147] ^ in[82]); 
    assign layer_0[1426] = in[181] ^ in[150]; 
    assign layer_0[1427] = in[210] | in[79]; 
    assign layer_0[1428] = ~(in[118] ^ in[132]); 
    assign layer_0[1429] = ~in[167]; 
    assign layer_0[1430] = ~(in[154] | in[171]); 
    assign layer_0[1431] = in[153]; 
    assign layer_0[1432] = in[111]; 
    assign layer_0[1433] = in[61] | in[57]; 
    assign layer_0[1434] = in[61] ^ in[27]; 
    assign layer_0[1435] = in[41]; 
    assign layer_0[1436] = in[245] & ~in[166]; 
    assign layer_0[1437] = ~(in[168] ^ in[234]); 
    assign layer_0[1438] = in[93] & ~in[30]; 
    assign layer_0[1439] = in[86]; 
    assign layer_0[1440] = ~(in[91] ^ in[89]); 
    assign layer_0[1441] = ~(in[116] ^ in[102]); 
    assign layer_0[1442] = ~(in[249] ^ in[246]); 
    assign layer_0[1443] = in[166] ^ in[243]; 
    assign layer_0[1444] = in[210] | in[7]; 
    assign layer_0[1445] = in[132] & ~in[119]; 
    assign layer_0[1446] = ~(in[116] ^ in[102]); 
    assign layer_0[1447] = ~(in[149] ^ in[147]); 
    assign layer_0[1448] = ~in[251]; 
    assign layer_0[1449] = ~(in[60] | in[127]); 
    assign layer_0[1450] = in[196] & ~in[215]; 
    assign layer_0[1451] = ~(in[12] ^ in[100]); 
    assign layer_0[1452] = in[165] | in[182]; 
    assign layer_0[1453] = in[169] ^ in[103]; 
    assign layer_0[1454] = ~in[89]; 
    assign layer_0[1455] = in[40] & ~in[163]; 
    assign layer_0[1456] = in[166] ^ in[227]; 
    assign layer_0[1457] = ~(in[105] ^ in[107]); 
    assign layer_0[1458] = ~(in[186] ^ in[189]); 
    assign layer_0[1459] = in[185] ^ in[213]; 
    assign layer_0[1460] = in[186] & ~in[137]; 
    assign layer_0[1461] = in[150]; 
    assign layer_0[1462] = ~(in[178] ^ in[121]); 
    assign layer_0[1463] = ~(in[195] | in[180]); 
    assign layer_0[1464] = ~in[150] | (in[150] & in[78]); 
    assign layer_0[1465] = ~in[133] | (in[133] & in[53]); 
    assign layer_0[1466] = ~(in[105] ^ in[137]); 
    assign layer_0[1467] = in[8] ^ in[55]; 
    assign layer_0[1468] = ~(in[154] ^ in[125]); 
    assign layer_0[1469] = in[104] & in[186]; 
    assign layer_0[1470] = in[88]; 
    assign layer_0[1471] = ~in[20] | (in[20] & in[83]); 
    assign layer_0[1472] = ~in[163] | (in[163] & in[79]); 
    assign layer_0[1473] = in[105] & ~in[135]; 
    assign layer_0[1474] = ~(in[123] ^ in[76]); 
    assign layer_0[1475] = in[30] | in[47]; 
    assign layer_0[1476] = in[8] | in[170]; 
    assign layer_0[1477] = in[9] | in[251]; 
    assign layer_0[1478] = ~(in[148] & in[167]); 
    assign layer_0[1479] = ~(in[6] | in[193]); 
    assign layer_0[1480] = ~(in[71] | in[93]); 
    assign layer_0[1481] = in[151] ^ in[197]; 
    assign layer_0[1482] = in[55] ^ in[215]; 
    assign layer_0[1483] = in[138] ^ in[156]; 
    assign layer_0[1484] = in[56] | in[110]; 
    assign layer_0[1485] = ~(in[196] ^ in[9]); 
    assign layer_0[1486] = in[26] | in[28]; 
    assign layer_0[1487] = ~(in[175] ^ in[206]); 
    assign layer_0[1488] = ~in[230] | (in[183] & in[230]); 
    assign layer_0[1489] = ~(in[233] | in[211]); 
    assign layer_0[1490] = ~(in[163] | in[148]); 
    assign layer_0[1491] = ~(in[218] ^ in[250]); 
    assign layer_0[1492] = ~(in[122] ^ in[155]); 
    assign layer_0[1493] = ~(in[235] ^ in[58]); 
    assign layer_0[1494] = in[108] & ~in[59]; 
    assign layer_0[1495] = ~in[110]; 
    assign layer_0[1496] = ~in[72] | (in[36] & in[72]); 
    assign layer_0[1497] = in[90] & ~in[61]; 
    assign layer_0[1498] = in[41] & ~in[151]; 
    assign layer_0[1499] = ~(in[164] | in[93]); 
    assign layer_0[1500] = in[102] | in[100]; 
    assign layer_0[1501] = in[107] & ~in[138]; 
    assign layer_0[1502] = ~(in[191] ^ in[179]); 
    assign layer_0[1503] = in[233]; 
    assign layer_0[1504] = ~(in[200] ^ in[53]); 
    assign layer_0[1505] = in[38] ^ in[69]; 
    assign layer_0[1506] = ~in[149] | (in[149] & in[132]); 
    assign layer_0[1507] = in[52] | in[74]; 
    assign layer_0[1508] = ~(in[86] ^ in[99]); 
    assign layer_0[1509] = in[47] | in[100]; 
    assign layer_0[1510] = in[198] ^ in[201]; 
    assign layer_0[1511] = ~(in[113] | in[101]); 
    assign layer_0[1512] = in[92] | in[238]; 
    assign layer_0[1513] = ~(in[177] | in[135]); 
    assign layer_0[1514] = in[86] | in[41]; 
    assign layer_0[1515] = ~(in[59] & in[245]); 
    assign layer_0[1516] = ~in[83]; 
    assign layer_0[1517] = ~(in[92] ^ in[171]); 
    assign layer_0[1518] = in[11]; 
    assign layer_0[1519] = in[147] ^ in[149]; 
    assign layer_0[1520] = ~(in[23] | in[61]); 
    assign layer_0[1521] = ~(in[31] ^ in[228]); 
    assign layer_0[1522] = ~(in[189] ^ in[156]); 
    assign layer_0[1523] = ~in[146]; 
    assign layer_0[1524] = ~in[247]; 
    assign layer_0[1525] = ~in[171]; 
    assign layer_0[1526] = in[67] | in[69]; 
    assign layer_0[1527] = in[93] ^ in[91]; 
    assign layer_0[1528] = ~in[122] | (in[122] & in[196]); 
    assign layer_0[1529] = in[200] & ~in[86]; 
    assign layer_0[1530] = in[152] | in[121]; 
    assign layer_0[1531] = ~in[194] | (in[196] & in[194]); 
    assign layer_0[1532] = in[73] & ~in[98]; 
    assign layer_0[1533] = in[150] ^ in[161]; 
    assign layer_0[1534] = in[146]; 
    assign layer_0[1535] = in[71] & ~in[42]; 
    assign layer_0[1536] = ~in[242] | (in[245] & in[242]); 
    assign layer_0[1537] = ~(in[70] ^ in[206]); 
    assign layer_0[1538] = ~in[126] | (in[126] & in[137]); 
    assign layer_0[1539] = in[165] | in[120]; 
    assign layer_0[1540] = in[117] ^ in[131]; 
    assign layer_0[1541] = ~(in[179] ^ in[237]); 
    assign layer_0[1542] = in[19] | in[65]; 
    assign layer_0[1543] = in[106] | in[147]; 
    assign layer_0[1544] = ~(in[72] & in[72]); 
    assign layer_0[1545] = ~(in[58] ^ in[89]); 
    assign layer_0[1546] = ~(in[93] & in[125]); 
    assign layer_0[1547] = in[140] & ~in[26]; 
    assign layer_0[1548] = in[78]; 
    assign layer_0[1549] = in[248] ^ in[228]; 
    assign layer_0[1550] = ~(in[170] | in[89]); 
    assign layer_0[1551] = ~in[114]; 
    assign layer_0[1552] = in[96] ^ in[190]; 
    assign layer_0[1553] = in[21] | in[9]; 
    assign layer_0[1554] = in[25] & ~in[57]; 
    assign layer_0[1555] = in[89]; 
    assign layer_0[1556] = in[196] | in[179]; 
    assign layer_0[1557] = in[60]; 
    assign layer_0[1558] = in[187]; 
    assign layer_0[1559] = in[115] ^ in[100]; 
    assign layer_0[1560] = ~in[153] | (in[141] & in[153]); 
    assign layer_0[1561] = ~in[9]; 
    assign layer_0[1562] = ~in[56]; 
    assign layer_0[1563] = in[61] & ~in[134]; 
    assign layer_0[1564] = in[216] & ~in[249]; 
    assign layer_0[1565] = ~(in[135] | in[148]); 
    assign layer_0[1566] = ~(in[30] | in[196]); 
    assign layer_0[1567] = in[211] ^ in[103]; 
    assign layer_0[1568] = ~(in[125] | in[114]); 
    assign layer_0[1569] = ~(in[129] | in[137]); 
    assign layer_0[1570] = in[55] & ~in[7]; 
    assign layer_0[1571] = ~in[40]; 
    assign layer_0[1572] = ~(in[38] ^ in[180]); 
    assign layer_0[1573] = ~(in[209] ^ in[133]); 
    assign layer_0[1574] = ~in[71] | (in[11] & in[71]); 
    assign layer_0[1575] = ~(in[83] ^ in[118]); 
    assign layer_0[1576] = in[245] ^ in[93]; 
    assign layer_0[1577] = ~(in[104] | in[211]); 
    assign layer_0[1578] = ~in[99] | (in[50] & in[99]); 
    assign layer_0[1579] = in[151] & ~in[61]; 
    assign layer_0[1580] = in[89] | in[76]; 
    assign layer_0[1581] = ~(in[73] | in[83]); 
    assign layer_0[1582] = ~(in[51] | in[94]); 
    assign layer_0[1583] = in[246]; 
    assign layer_0[1584] = ~(in[8] | in[20]); 
    assign layer_0[1585] = ~in[138] | (in[119] & in[138]); 
    assign layer_0[1586] = ~(in[151] | in[135]); 
    assign layer_0[1587] = ~(in[219] & in[73]); 
    assign layer_0[1588] = in[164]; 
    assign layer_0[1589] = in[101] | in[242]; 
    assign layer_0[1590] = ~in[137] | (in[22] & in[137]); 
    assign layer_0[1591] = ~in[44]; 
    assign layer_0[1592] = ~(in[232] ^ in[249]); 
    assign layer_0[1593] = ~in[88] | (in[88] & in[12]); 
    assign layer_0[1594] = in[121] ^ in[168]; 
    assign layer_0[1595] = in[119] | in[108]; 
    assign layer_0[1596] = in[152]; 
    assign layer_0[1597] = in[229] | in[214]; 
    assign layer_0[1598] = in[74] & ~in[114]; 
    assign layer_0[1599] = in[120] & ~in[140]; 
    assign layer_0[1600] = ~(in[41] | in[61]); 
    assign layer_0[1601] = ~(in[51] ^ in[22]); 
    assign layer_0[1602] = ~in[194]; 
    assign layer_0[1603] = in[118] | in[86]; 
    assign layer_0[1604] = ~(in[26] | in[45]); 
    assign layer_0[1605] = ~(in[86] ^ in[98]); 
    assign layer_0[1606] = in[137] & ~in[139]; 
    assign layer_0[1607] = ~in[87] | (in[118] & in[87]); 
    assign layer_0[1608] = ~(in[218] | in[46]); 
    assign layer_0[1609] = ~in[187] | (in[187] & in[210]); 
    assign layer_0[1610] = in[101] | in[20]; 
    assign layer_0[1611] = in[130] | in[115]; 
    assign layer_0[1612] = in[149] ^ in[118]; 
    assign layer_0[1613] = in[76] | in[251]; 
    assign layer_0[1614] = in[137] ^ in[35]; 
    assign layer_0[1615] = ~in[115] | (in[115] & in[80]); 
    assign layer_0[1616] = in[151]; 
    assign layer_0[1617] = in[120] ^ in[67]; 
    assign layer_0[1618] = in[89] | in[94]; 
    assign layer_0[1619] = in[228] ^ in[182]; 
    assign layer_0[1620] = in[185] | in[227]; 
    assign layer_0[1621] = ~(in[91] ^ in[93]); 
    assign layer_0[1622] = in[42] ^ in[75]; 
    assign layer_0[1623] = in[231] | in[106]; 
    assign layer_0[1624] = in[215] & ~in[228]; 
    assign layer_0[1625] = ~in[213] | (in[9] & in[213]); 
    assign layer_0[1626] = in[89] & ~in[76]; 
    assign layer_0[1627] = in[205] ^ in[173]; 
    assign layer_0[1628] = in[169] & ~in[211]; 
    assign layer_0[1629] = in[230] ^ in[135]; 
    assign layer_0[1630] = ~(in[37] ^ in[67]); 
    assign layer_0[1631] = ~in[59] | (in[59] & in[85]); 
    assign layer_0[1632] = in[113] ^ in[102]; 
    assign layer_0[1633] = in[237] | in[133]; 
    assign layer_0[1634] = ~(in[241] | in[100]); 
    assign layer_0[1635] = in[115] & ~in[193]; 
    assign layer_0[1636] = ~in[219]; 
    assign layer_0[1637] = ~(in[142] | in[74]); 
    assign layer_0[1638] = in[249] ^ in[217]; 
    assign layer_0[1639] = in[101] ^ in[99]; 
    assign layer_0[1640] = ~(in[78] ^ in[74]); 
    assign layer_0[1641] = in[111] | in[126]; 
    assign layer_0[1642] = ~(in[135] ^ in[104]); 
    assign layer_0[1643] = ~(in[248] ^ in[185]); 
    assign layer_0[1644] = ~(in[126] | in[198]); 
    assign layer_0[1645] = ~(in[53] & in[235]); 
    assign layer_0[1646] = in[88]; 
    assign layer_0[1647] = in[98] | in[169]; 
    assign layer_0[1648] = in[53]; 
    assign layer_0[1649] = ~in[122] | (in[122] & in[28]); 
    assign layer_0[1650] = in[114] ^ in[116]; 
    assign layer_0[1651] = ~(in[141] ^ in[143]); 
    assign layer_0[1652] = in[171] ^ in[242]; 
    assign layer_0[1653] = in[197] & ~in[110]; 
    assign layer_0[1654] = in[126] ^ in[12]; 
    assign layer_0[1655] = ~in[6]; 
    assign layer_0[1656] = ~in[90]; 
    assign layer_0[1657] = ~(in[140] | in[122]); 
    assign layer_0[1658] = ~(in[115] ^ in[117]); 
    assign layer_0[1659] = in[20] ^ in[196]; 
    assign layer_0[1660] = in[104] ^ in[55]; 
    assign layer_0[1661] = ~(in[11] ^ in[119]); 
    assign layer_0[1662] = ~(in[8] ^ in[29]); 
    assign layer_0[1663] = in[106] ^ in[108]; 
    assign layer_0[1664] = in[132] | in[101]; 
    assign layer_0[1665] = ~(in[53] ^ in[180]); 
    assign layer_0[1666] = ~(in[116] | in[108]); 
    assign layer_0[1667] = ~in[152] | (in[152] & in[7]); 
    assign layer_0[1668] = in[11]; 
    assign layer_0[1669] = ~(in[147] ^ in[165]); 
    assign layer_0[1670] = ~(in[43] ^ in[75]); 
    assign layer_0[1671] = ~(in[62] ^ in[27]); 
    assign layer_0[1672] = ~in[57] | (in[57] & in[167]); 
    assign layer_0[1673] = in[121] | in[30]; 
    assign layer_0[1674] = ~(in[58] ^ in[89]); 
    assign layer_0[1675] = in[137] & ~in[234]; 
    assign layer_0[1676] = in[25] | in[221]; 
    assign layer_0[1677] = ~(in[117] | in[47]); 
    assign layer_0[1678] = in[194] ^ in[60]; 
    assign layer_0[1679] = in[211] ^ in[226]; 
    assign layer_0[1680] = in[98]; 
    assign layer_0[1681] = in[153] ^ in[122]; 
    assign layer_0[1682] = ~in[124]; 
    assign layer_0[1683] = in[183] ^ in[180]; 
    assign layer_0[1684] = ~(in[10] | in[41]); 
    assign layer_0[1685] = in[130]; 
    assign layer_0[1686] = ~in[185]; 
    assign layer_0[1687] = in[58] ^ in[234]; 
    assign layer_0[1688] = in[164] | in[204]; 
    assign layer_0[1689] = ~in[105]; 
    assign layer_0[1690] = ~(in[134] ^ in[200]); 
    assign layer_0[1691] = ~(in[54] ^ in[38]); 
    assign layer_0[1692] = in[107] ^ in[82]; 
    assign layer_0[1693] = in[150] ^ in[116]; 
    assign layer_0[1694] = ~(in[94] | in[90]); 
    assign layer_0[1695] = ~in[57] | (in[57] & in[155]); 
    assign layer_0[1696] = ~in[201] | (in[201] & in[213]); 
    assign layer_0[1697] = ~(in[170] ^ in[73]); 
    assign layer_0[1698] = in[56]; 
    assign layer_0[1699] = in[113] | in[72]; 
    assign layer_0[1700] = in[154] | in[186]; 
    assign layer_0[1701] = in[139] & ~in[196]; 
    assign layer_0[1702] = in[139] ^ in[73]; 
    assign layer_0[1703] = in[69] ^ in[73]; 
    assign layer_0[1704] = in[61] & ~in[139]; 
    assign layer_0[1705] = in[130]; 
    assign layer_0[1706] = in[123] ^ in[49]; 
    assign layer_0[1707] = in[147] & ~in[229]; 
    assign layer_0[1708] = ~(in[221] | in[78]); 
    assign layer_0[1709] = in[23] ^ in[219]; 
    assign layer_0[1710] = ~in[88]; 
    assign layer_0[1711] = ~(in[177] ^ in[225]); 
    assign layer_0[1712] = ~(in[185] ^ in[182]); 
    assign layer_0[1713] = ~(in[69] ^ in[185]); 
    assign layer_0[1714] = in[77] ^ in[75]; 
    assign layer_0[1715] = ~in[139]; 
    assign layer_0[1716] = ~in[231] | (in[231] & in[181]); 
    assign layer_0[1717] = ~(in[168] & in[232]); 
    assign layer_0[1718] = ~(in[51] ^ in[75]); 
    assign layer_0[1719] = in[130] & ~in[65]; 
    assign layer_0[1720] = in[163] | in[166]; 
    assign layer_0[1721] = ~(in[167] | in[211]); 
    assign layer_0[1722] = ~in[158]; 
    assign layer_0[1723] = in[55] | in[102]; 
    assign layer_0[1724] = ~(in[251] | in[152]); 
    assign layer_0[1725] = ~(in[83] ^ in[69]); 
    assign layer_0[1726] = ~in[216] | (in[141] & in[216]); 
    assign layer_0[1727] = in[82] | in[182]; 
    assign layer_0[1728] = in[141] ^ in[147]; 
    assign layer_0[1729] = in[211] & in[164]; 
    assign layer_0[1730] = in[198] | in[167]; 
    assign layer_0[1731] = ~(in[36] ^ in[85]); 
    assign layer_0[1732] = in[162] | in[85]; 
    assign layer_0[1733] = ~(in[13] | in[231]); 
    assign layer_0[1734] = in[58] ^ in[121]; 
    assign layer_0[1735] = in[25]; 
    assign layer_0[1736] = ~(in[36] ^ in[25]); 
    assign layer_0[1737] = ~(in[155] | in[53]); 
    assign layer_0[1738] = in[145] ^ in[6]; 
    assign layer_0[1739] = ~(in[247] | in[231]); 
    assign layer_0[1740] = in[9]; 
    assign layer_0[1741] = ~in[123] | (in[123] & in[167]); 
    assign layer_0[1742] = in[44] ^ in[57]; 
    assign layer_0[1743] = ~(in[152] | in[150]); 
    assign layer_0[1744] = in[181] ^ in[183]; 
    assign layer_0[1745] = in[164] & in[132]; 
    assign layer_0[1746] = ~(in[116] ^ in[20]); 
    assign layer_0[1747] = in[93] | in[72]; 
    assign layer_0[1748] = ~in[165] | (in[245] & in[165]); 
    assign layer_0[1749] = ~(in[200] ^ in[243]); 
    assign layer_0[1750] = ~in[68]; 
    assign layer_0[1751] = in[148] | in[228]; 
    assign layer_0[1752] = in[90] & in[148]; 
    assign layer_0[1753] = in[38] ^ in[69]; 
    assign layer_0[1754] = ~in[138] | (in[138] & in[197]); 
    assign layer_0[1755] = ~(in[213] ^ in[243]); 
    assign layer_0[1756] = ~(in[165] ^ in[163]); 
    assign layer_0[1757] = ~(in[126] | in[111]); 
    assign layer_0[1758] = in[183] ^ in[180]; 
    assign layer_0[1759] = in[206] | in[72]; 
    assign layer_0[1760] = ~in[193]; 
    assign layer_0[1761] = ~(in[21] | in[11]); 
    assign layer_0[1762] = ~(in[102] & in[151]); 
    assign layer_0[1763] = in[116] & ~in[181]; 
    assign layer_0[1764] = in[87] ^ in[55]; 
    assign layer_0[1765] = ~in[89] | (in[89] & in[180]); 
    assign layer_0[1766] = in[189] ^ in[41]; 
    assign layer_0[1767] = ~(in[229] | in[140]); 
    assign layer_0[1768] = ~(in[181] ^ in[85]); 
    assign layer_0[1769] = in[9]; 
    assign layer_0[1770] = ~in[132]; 
    assign layer_0[1771] = in[70] | in[98]; 
    assign layer_0[1772] = ~(in[208] ^ in[5]); 
    assign layer_0[1773] = in[90] ^ in[138]; 
    assign layer_0[1774] = in[158] | in[241]; 
    assign layer_0[1775] = ~(in[194] | in[101]); 
    assign layer_0[1776] = ~in[70]; 
    assign layer_0[1777] = ~in[133] | (in[133] & in[151]); 
    assign layer_0[1778] = ~in[167]; 
    assign layer_0[1779] = ~in[175]; 
    assign layer_0[1780] = in[119] & ~in[56]; 
    assign layer_0[1781] = in[78] ^ in[57]; 
    assign layer_0[1782] = ~(in[106] ^ in[93]); 
    assign layer_0[1783] = ~in[211]; 
    assign layer_0[1784] = in[173] ^ in[139]; 
    assign layer_0[1785] = in[204] ^ in[201]; 
    assign layer_0[1786] = in[141] | in[225]; 
    assign layer_0[1787] = in[230] ^ in[88]; 
    assign layer_0[1788] = ~(in[194] ^ in[221]); 
    assign layer_0[1789] = ~(in[170] ^ in[203]); 
    assign layer_0[1790] = ~(in[153] | in[184]); 
    assign layer_0[1791] = in[36] | in[91]; 
    assign layer_0[1792] = ~(in[198] ^ in[154]); 
    assign layer_0[1793] = in[88] ^ in[232]; 
    assign layer_0[1794] = ~(in[179] | in[214]); 
    assign layer_0[1795] = ~(in[6] | in[155]); 
    assign layer_0[1796] = ~(in[179] | in[57]); 
    assign layer_0[1797] = ~(in[99] ^ in[53]); 
    assign layer_0[1798] = ~(in[156] | in[92]); 
    assign layer_0[1799] = ~(in[155] ^ in[46]); 
    assign layer_0[1800] = in[101]; 
    assign layer_0[1801] = ~in[55] | (in[55] & in[199]); 
    assign layer_0[1802] = ~(in[214] | in[131]); 
    assign layer_0[1803] = ~(in[118] | in[133]); 
    assign layer_0[1804] = in[116] & ~in[164]; 
    assign layer_0[1805] = ~(in[214] ^ in[245]); 
    assign layer_0[1806] = in[122] ^ in[166]; 
    assign layer_0[1807] = ~in[215]; 
    assign layer_0[1808] = in[161]; 
    assign layer_0[1809] = in[103] ^ in[73]; 
    assign layer_0[1810] = ~(in[162] | in[178]); 
    assign layer_0[1811] = ~(in[186] | in[101]); 
    assign layer_0[1812] = ~(in[98] | in[242]); 
    assign layer_0[1813] = ~in[170] | (in[170] & in[53]); 
    assign layer_0[1814] = ~(in[183] ^ in[21]); 
    assign layer_0[1815] = ~in[73] | (in[11] & in[73]); 
    assign layer_0[1816] = ~(in[122] & in[120]); 
    assign layer_0[1817] = ~in[90] | (in[90] & in[193]); 
    assign layer_0[1818] = in[100] | in[139]; 
    assign layer_0[1819] = in[24] ^ in[70]; 
    assign layer_0[1820] = in[136] & ~in[125]; 
    assign layer_0[1821] = in[201] ^ in[170]; 
    assign layer_0[1822] = in[148] | in[183]; 
    assign layer_0[1823] = ~in[103]; 
    assign layer_0[1824] = in[139] ^ in[77]; 
    assign layer_0[1825] = ~in[29] | (in[133] & in[29]); 
    assign layer_0[1826] = ~in[151] | (in[179] & in[151]); 
    assign layer_0[1827] = in[11] | in[223]; 
    assign layer_0[1828] = ~in[151] | (in[151] & in[74]); 
    assign layer_0[1829] = in[78] ^ in[250]; 
    assign layer_0[1830] = ~(in[117] ^ in[121]); 
    assign layer_0[1831] = ~(in[235] ^ in[60]); 
    assign layer_0[1832] = ~(in[218] | in[177]); 
    assign layer_0[1833] = ~(in[134] | in[116]); 
    assign layer_0[1834] = ~(in[113] ^ in[103]); 
    assign layer_0[1835] = in[59] & ~in[118]; 
    assign layer_0[1836] = ~(in[157] | in[71]); 
    assign layer_0[1837] = in[93] & in[179]; 
    assign layer_0[1838] = ~(in[153] ^ in[82]); 
    assign layer_0[1839] = ~in[244]; 
    assign layer_0[1840] = ~(in[41] | in[43]); 
    assign layer_0[1841] = in[213] & ~in[122]; 
    assign layer_0[1842] = ~(in[119] | in[28]); 
    assign layer_0[1843] = ~(in[89] ^ in[58]); 
    assign layer_0[1844] = in[66] | in[35]; 
    assign layer_0[1845] = ~(in[198] ^ in[248]); 
    assign layer_0[1846] = ~(in[140] | in[109]); 
    assign layer_0[1847] = ~(in[244] ^ in[252]); 
    assign layer_0[1848] = in[79] ^ in[248]; 
    assign layer_0[1849] = ~(in[188] | in[185]); 
    assign layer_0[1850] = ~in[124]; 
    assign layer_0[1851] = ~(in[118] | in[149]); 
    assign layer_0[1852] = in[90] & ~in[26]; 
    assign layer_0[1853] = ~(in[163] ^ in[123]); 
    assign layer_0[1854] = in[212] ^ in[198]; 
    assign layer_0[1855] = ~in[153]; 
    assign layer_0[1856] = ~in[122] | (in[93] & in[122]); 
    assign layer_0[1857] = ~(in[69] | in[86]); 
    assign layer_0[1858] = ~in[23] | (in[23] & in[87]); 
    assign layer_0[1859] = ~in[217] | (in[198] & in[217]); 
    assign layer_0[1860] = in[72] | in[74]; 
    assign layer_0[1861] = in[166]; 
    assign layer_0[1862] = in[211] & ~in[88]; 
    assign layer_0[1863] = ~(in[204] ^ in[235]); 
    assign layer_0[1864] = ~(in[53] | in[91]); 
    assign layer_0[1865] = ~(in[151] ^ in[120]); 
    assign layer_0[1866] = ~in[20] | (in[20] & in[181]); 
    assign layer_0[1867] = in[137] | in[252]; 
    assign layer_0[1868] = in[182] ^ in[228]; 
    assign layer_0[1869] = in[158] ^ in[215]; 
    assign layer_0[1870] = ~(in[120] ^ in[211]); 
    assign layer_0[1871] = ~(in[165] ^ in[130]); 
    assign layer_0[1872] = ~in[233] | (in[233] & in[125]); 
    assign layer_0[1873] = ~(in[164] ^ in[229]); 
    assign layer_0[1874] = in[47] & ~in[140]; 
    assign layer_0[1875] = ~(in[36] | in[67]); 
    assign layer_0[1876] = in[227] ^ in[243]; 
    assign layer_0[1877] = ~(in[188] | in[203]); 
    assign layer_0[1878] = in[88] & ~in[213]; 
    assign layer_0[1879] = in[221] ^ in[194]; 
    assign layer_0[1880] = ~(in[54] ^ in[99]); 
    assign layer_0[1881] = in[244] | in[237]; 
    assign layer_0[1882] = ~in[202]; 
    assign layer_0[1883] = in[146] ^ in[148]; 
    assign layer_0[1884] = in[88]; 
    assign layer_0[1885] = ~(in[146] | in[201]); 
    assign layer_0[1886] = in[110] & ~in[242]; 
    assign layer_0[1887] = ~(in[246] ^ in[188]); 
    assign layer_0[1888] = ~(in[227] ^ in[24]); 
    assign layer_0[1889] = ~in[5]; 
    assign layer_0[1890] = ~(in[106] ^ in[124]); 
    assign layer_0[1891] = ~in[135] | (in[135] & in[141]); 
    assign layer_0[1892] = ~(in[143] ^ in[40]); 
    assign layer_0[1893] = in[35] | in[6]; 
    assign layer_0[1894] = in[24]; 
    assign layer_0[1895] = ~(in[131] ^ in[119]); 
    assign layer_0[1896] = ~(in[205] ^ in[162]); 
    assign layer_0[1897] = ~in[200] | (in[57] & in[200]); 
    assign layer_0[1898] = in[195] & ~in[188]; 
    assign layer_0[1899] = ~(in[228] ^ in[197]); 
    assign layer_0[1900] = in[247] ^ in[196]; 
    assign layer_0[1901] = in[247] ^ in[26]; 
    assign layer_0[1902] = ~(in[135] ^ in[40]); 
    assign layer_0[1903] = in[93] | in[61]; 
    assign layer_0[1904] = ~(in[63] ^ in[46]); 
    assign layer_0[1905] = ~in[187]; 
    assign layer_0[1906] = ~(in[216] | in[249]); 
    assign layer_0[1907] = ~in[234] | (in[85] & in[234]); 
    assign layer_0[1908] = in[60] ^ in[249]; 
    assign layer_0[1909] = in[163] | in[196]; 
    assign layer_0[1910] = ~(in[182] ^ in[163]); 
    assign layer_0[1911] = ~in[120]; 
    assign layer_0[1912] = ~in[183] | (in[183] & in[249]); 
    assign layer_0[1913] = in[211] ^ in[233]; 
    assign layer_0[1914] = in[144] | in[194]; 
    assign layer_0[1915] = ~in[137] | (in[137] & in[218]); 
    assign layer_0[1916] = ~(in[156] ^ in[122]); 
    assign layer_0[1917] = ~in[137]; 
    assign layer_0[1918] = ~(in[117] ^ in[102]); 
    assign layer_0[1919] = ~in[152]; 
    assign layer_0[1920] = ~(in[101] ^ in[180]); 
    assign layer_0[1921] = ~(in[85] ^ in[199]); 
    assign layer_0[1922] = ~in[202] | (in[133] & in[202]); 
    assign layer_0[1923] = in[174] ^ in[118]; 
    assign layer_0[1924] = ~(in[196] | in[231]); 
    assign layer_0[1925] = ~in[71]; 
    assign layer_0[1926] = ~(in[86] ^ in[157]); 
    assign layer_0[1927] = in[244] ^ in[129]; 
    assign layer_0[1928] = ~in[72]; 
    assign layer_0[1929] = ~(in[116] ^ in[165]); 
    assign layer_0[1930] = in[74] & ~in[136]; 
    assign layer_0[1931] = ~(in[166] | in[45]); 
    assign layer_0[1932] = in[153]; 
    assign layer_0[1933] = ~in[201]; 
    assign layer_0[1934] = ~in[89] | (in[89] & in[106]); 
    assign layer_0[1935] = ~in[138]; 
    assign layer_0[1936] = in[117] ^ in[103]; 
    assign layer_0[1937] = ~(in[207] ^ in[29]); 
    assign layer_0[1938] = ~(in[187] ^ in[209]); 
    assign layer_0[1939] = ~in[134] | (in[134] & in[140]); 
    assign layer_0[1940] = in[226] ^ in[244]; 
    assign layer_0[1941] = in[146] | in[92]; 
    assign layer_0[1942] = in[94] ^ in[92]; 
    assign layer_0[1943] = in[88] ^ in[73]; 
    assign layer_0[1944] = ~(in[95] | in[79]); 
    assign layer_0[1945] = in[156]; 
    assign layer_0[1946] = ~in[22] | (in[99] & in[22]); 
    assign layer_0[1947] = ~(in[165] ^ in[162]); 
    assign layer_0[1948] = in[55] ^ in[100]; 
    assign layer_0[1949] = ~(in[214] ^ in[6]); 
    assign layer_0[1950] = in[68] | in[41]; 
    assign layer_0[1951] = in[198] ^ in[244]; 
    assign layer_0[1952] = ~(in[106] ^ in[137]); 
    assign layer_0[1953] = ~in[143]; 
    assign layer_0[1954] = ~(in[172] | in[201]); 
    assign layer_0[1955] = in[50] ^ in[20]; 
    assign layer_0[1956] = ~(in[94] ^ in[107]); 
    assign layer_0[1957] = ~(in[139] | in[101]); 
    assign layer_0[1958] = ~(in[28] | in[94]); 
    assign layer_0[1959] = ~(in[166] ^ in[164]); 
    assign layer_0[1960] = ~in[60] | (in[226] & in[60]); 
    assign layer_0[1961] = in[153] & ~in[232]; 
    assign layer_0[1962] = in[72] & in[75]; 
    assign layer_0[1963] = in[95] ^ in[92]; 
    assign layer_0[1964] = in[88] ^ in[102]; 
    assign layer_0[1965] = ~(in[129] ^ in[168]); 
    assign layer_0[1966] = in[231]; 
    assign layer_0[1967] = in[60] ^ in[54]; 
    assign layer_0[1968] = in[102]; 
    assign layer_0[1969] = in[149]; 
    assign layer_0[1970] = in[152] ^ in[105]; 
    assign layer_0[1971] = ~(in[110] | in[124]); 
    assign layer_0[1972] = in[60] & in[213]; 
    assign layer_0[1973] = ~(in[198] | in[193]); 
    assign layer_0[1974] = in[139] | in[78]; 
    assign layer_0[1975] = in[195] ^ in[178]; 
    assign layer_0[1976] = in[79]; 
    assign layer_0[1977] = in[73] & ~in[23]; 
    assign layer_0[1978] = in[86] & ~in[37]; 
    assign layer_0[1979] = ~(in[28] ^ in[73]); 
    assign layer_0[1980] = ~in[34]; 
    assign layer_0[1981] = ~(in[24] ^ in[71]); 
    assign layer_0[1982] = ~(in[146] ^ in[148]); 
    assign layer_0[1983] = in[162] ^ in[164]; 
    assign layer_0[1984] = ~(in[232] ^ in[108]); 
    assign layer_0[1985] = in[189] | in[56]; 
    assign layer_0[1986] = in[202] ^ in[154]; 
    assign layer_0[1987] = in[138] & ~in[132]; 
    assign layer_0[1988] = in[76] ^ in[51]; 
    assign layer_0[1989] = ~(in[141] ^ in[171]); 
    assign layer_0[1990] = in[72] & ~in[151]; 
    assign layer_0[1991] = in[103] ^ in[185]; 
    assign layer_0[1992] = ~(in[250] ^ in[206]); 
    assign layer_0[1993] = ~(in[163] ^ in[133]); 
    assign layer_0[1994] = in[11]; 
    assign layer_0[1995] = ~in[199] | (in[199] & in[197]); 
    assign layer_0[1996] = ~(in[67] | in[87]); 
    assign layer_0[1997] = in[75] ^ in[77]; 
    assign layer_0[1998] = in[28] | in[179]; 
    assign layer_0[1999] = ~(in[65] ^ in[212]); 
    assign layer_0[2000] = ~in[70] | (in[136] & in[70]); 
    assign layer_0[2001] = ~in[85]; 
    assign layer_0[2002] = in[170] ^ in[26]; 
    assign layer_0[2003] = in[131] | in[27]; 
    assign layer_0[2004] = ~in[8] | (in[41] & in[8]); 
    assign layer_0[2005] = in[170]; 
    assign layer_0[2006] = in[171] | in[46]; 
    assign layer_0[2007] = in[169] ^ in[138]; 
    assign layer_0[2008] = in[70] ^ in[39]; 
    assign layer_0[2009] = in[58] ^ in[88]; 
    assign layer_0[2010] = ~in[178]; 
    assign layer_0[2011] = in[38] & ~in[168]; 
    assign layer_0[2012] = ~in[212]; 
    assign layer_0[2013] = in[166] ^ in[211]; 
    assign layer_0[2014] = in[198]; 
    assign layer_0[2015] = in[26] ^ in[45]; 
    assign layer_0[2016] = in[38] & ~in[74]; 
    assign layer_0[2017] = ~(in[217] ^ in[214]); 
    assign layer_0[2018] = in[123] ^ in[37]; 
    assign layer_0[2019] = ~(in[71] ^ in[213]); 
    assign layer_0[2020] = ~(in[121] ^ in[146]); 
    assign layer_0[2021] = in[83] & ~in[199]; 
    assign layer_0[2022] = ~in[143]; 
    assign layer_0[2023] = in[244] & ~in[180]; 
    assign layer_0[2024] = in[115]; 
    assign layer_0[2025] = in[124] | in[99]; 
    assign layer_0[2026] = in[99] ^ in[78]; 
    assign layer_0[2027] = ~in[132] | (in[120] & in[132]); 
    assign layer_0[2028] = ~in[122] | (in[122] & in[41]); 
    assign layer_0[2029] = in[134] & ~in[132]; 
    assign layer_0[2030] = in[25] ^ in[127]; 
    assign layer_0[2031] = in[214] | in[229]; 
    assign layer_0[2032] = ~(in[181] ^ in[164]); 
    assign layer_0[2033] = in[10]; 
    assign layer_0[2034] = ~(in[165] ^ in[162]); 
    assign layer_0[2035] = in[184]; 
    assign layer_0[2036] = ~(in[171] | in[188]); 
    assign layer_0[2037] = in[184] & ~in[134]; 
    assign layer_0[2038] = ~(in[251] ^ in[181]); 
    assign layer_0[2039] = in[249] ^ in[217]; 
    assign layer_0[2040] = in[253] | in[113]; 
    assign layer_0[2041] = in[165] ^ in[147]; 
    assign layer_0[2042] = ~(in[29] ^ in[11]); 
    assign layer_0[2043] = ~(in[213] ^ in[202]); 
    assign layer_0[2044] = ~(in[173] ^ in[230]); 
    assign layer_0[2045] = in[184] & ~in[212]; 
    assign layer_0[2046] = ~in[220]; 
    assign layer_0[2047] = ~(in[26] ^ in[184]); 
    assign layer_0[2048] = ~(in[23] | in[219]); 
    assign layer_0[2049] = ~(in[75] ^ in[87]); 
    assign layer_0[2050] = ~(in[28] | in[8]); 
    assign layer_0[2051] = in[90] & ~in[211]; 
    assign layer_0[2052] = in[54]; 
    assign layer_0[2053] = in[126] | in[228]; 
    assign layer_0[2054] = ~(in[244] | in[249]); 
    assign layer_0[2055] = in[100] & ~in[118]; 
    assign layer_0[2056] = ~(in[232] ^ in[201]); 
    assign layer_0[2057] = ~(in[210] | in[251]); 
    assign layer_0[2058] = ~(in[57] ^ in[27]); 
    assign layer_0[2059] = in[30] | in[236]; 
    assign layer_0[2060] = in[150] | in[26]; 
    assign layer_0[2061] = in[190]; 
    assign layer_0[2062] = in[108] & ~in[215]; 
    assign layer_0[2063] = in[114] ^ in[57]; 
    assign layer_0[2064] = ~in[105] | (in[105] & in[151]); 
    assign layer_0[2065] = ~(in[248] | in[63]); 
    assign layer_0[2066] = ~in[21] | (in[21] & in[203]); 
    assign layer_0[2067] = in[245]; 
    assign layer_0[2068] = in[120] ^ in[86]; 
    assign layer_0[2069] = in[25] | in[38]; 
    assign layer_0[2070] = in[222] ^ in[191]; 
    assign layer_0[2071] = in[176] | in[243]; 
    assign layer_0[2072] = in[50] | in[139]; 
    assign layer_0[2073] = in[119] ^ in[150]; 
    assign layer_0[2074] = in[149] ^ in[107]; 
    assign layer_0[2075] = in[163] & in[204]; 
    assign layer_0[2076] = ~(in[121] ^ in[146]); 
    assign layer_0[2077] = in[104] & ~in[158]; 
    assign layer_0[2078] = in[245] | in[120]; 
    assign layer_0[2079] = ~(in[154] | in[21]); 
    assign layer_0[2080] = in[52] | in[34]; 
    assign layer_0[2081] = ~(in[52] ^ in[81]); 
    assign layer_0[2082] = ~(in[98] | in[116]); 
    assign layer_0[2083] = ~in[234]; 
    assign layer_0[2084] = ~(in[235] ^ in[205]); 
    assign layer_0[2085] = in[102] & ~in[148]; 
    assign layer_0[2086] = in[185] | in[109]; 
    assign layer_0[2087] = ~in[88] | (in[88] & in[60]); 
    assign layer_0[2088] = ~in[51]; 
    assign layer_0[2089] = in[85] ^ in[98]; 
    assign layer_0[2090] = in[25] | in[88]; 
    assign layer_0[2091] = in[91] & ~in[26]; 
    assign layer_0[2092] = ~(in[135] ^ in[152]); 
    assign layer_0[2093] = ~(in[132] | in[142]); 
    assign layer_0[2094] = ~(in[219] ^ in[251]); 
    assign layer_0[2095] = in[250] | in[51]; 
    assign layer_0[2096] = in[116] | in[189]; 
    assign layer_0[2097] = in[143] & ~in[120]; 
    assign layer_0[2098] = ~(in[182] | in[180]); 
    assign layer_0[2099] = ~in[52] | (in[39] & in[52]); 
    assign layer_0[2100] = ~in[197] | (in[197] & in[84]); 
    assign layer_0[2101] = ~in[57] | (in[187] & in[57]); 
    assign layer_0[2102] = ~(in[180] ^ in[149]); 
    assign layer_0[2103] = in[199] & ~in[46]; 
    assign layer_0[2104] = in[235] ^ in[59]; 
    assign layer_0[2105] = ~(in[219] ^ in[249]); 
    assign layer_0[2106] = ~in[135] | (in[135] & in[117]); 
    assign layer_0[2107] = ~(in[248] | in[249]); 
    assign layer_0[2108] = ~in[185]; 
    assign layer_0[2109] = in[125]; 
    assign layer_0[2110] = ~(in[102] | in[101]); 
    assign layer_0[2111] = ~(in[248] ^ in[59]); 
    assign layer_0[2112] = in[105] & ~in[70]; 
    assign layer_0[2113] = ~in[98] | (in[98] & in[137]); 
    assign layer_0[2114] = ~in[203] | (in[203] & in[82]); 
    assign layer_0[2115] = in[114] | in[91]; 
    assign layer_0[2116] = ~(in[150] ^ in[132]); 
    assign layer_0[2117] = in[72] & ~in[23]; 
    assign layer_0[2118] = in[73] ^ in[97]; 
    assign layer_0[2119] = ~(in[217] ^ in[76]); 
    assign layer_0[2120] = in[242] ^ in[212]; 
    assign layer_0[2121] = ~(in[207] ^ in[226]); 
    assign layer_0[2122] = in[150] & ~in[177]; 
    assign layer_0[2123] = in[108] | in[142]; 
    assign layer_0[2124] = in[154] ^ in[122]; 
    assign layer_0[2125] = in[79] ^ in[36]; 
    assign layer_0[2126] = in[116] & ~in[91]; 
    assign layer_0[2127] = ~(in[120] ^ in[151]); 
    assign layer_0[2128] = in[183] ^ in[100]; 
    assign layer_0[2129] = ~(in[199] ^ in[247]); 
    assign layer_0[2130] = ~in[166]; 
    assign layer_0[2131] = ~in[119]; 
    assign layer_0[2132] = ~in[5]; 
    assign layer_0[2133] = in[107] ^ in[110]; 
    assign layer_0[2134] = in[184] ^ in[119]; 
    assign layer_0[2135] = in[150]; 
    assign layer_0[2136] = in[152] & ~in[63]; 
    assign layer_0[2137] = in[185] | in[30]; 
    assign layer_0[2138] = ~(in[200] ^ in[88]); 
    assign layer_0[2139] = in[139] ^ in[104]; 
    assign layer_0[2140] = in[61]; 
    assign layer_0[2141] = ~(in[54] ^ in[23]); 
    assign layer_0[2142] = ~in[179] | (in[149] & in[179]); 
    assign layer_0[2143] = in[40] | in[72]; 
    assign layer_0[2144] = in[184]; 
    assign layer_0[2145] = in[137]; 
    assign layer_0[2146] = in[21] ^ in[60]; 
    assign layer_0[2147] = in[244] ^ in[151]; 
    assign layer_0[2148] = in[178] | in[167]; 
    assign layer_0[2149] = in[76] ^ in[74]; 
    assign layer_0[2150] = in[152] ^ in[199]; 
    assign layer_0[2151] = in[250] ^ in[76]; 
    assign layer_0[2152] = in[137] | in[139]; 
    assign layer_0[2153] = in[58] & ~in[52]; 
    assign layer_0[2154] = in[222] | in[194]; 
    assign layer_0[2155] = in[167] & ~in[247]; 
    assign layer_0[2156] = ~in[120] | (in[41] & in[120]); 
    assign layer_0[2157] = ~(in[169] | in[105]); 
    assign layer_0[2158] = in[233] ^ in[197]; 
    assign layer_0[2159] = ~in[165]; 
    assign layer_0[2160] = ~(in[212] | in[109]); 
    assign layer_0[2161] = in[119] & ~in[69]; 
    assign layer_0[2162] = in[90] & ~in[233]; 
    assign layer_0[2163] = in[100] & ~in[119]; 
    assign layer_0[2164] = ~(in[230] ^ in[248]); 
    assign layer_0[2165] = in[203] & ~in[81]; 
    assign layer_0[2166] = ~(in[90] ^ in[106]); 
    assign layer_0[2167] = in[76] & ~in[166]; 
    assign layer_0[2168] = ~(in[127] ^ in[150]); 
    assign layer_0[2169] = in[133] | in[42]; 
    assign layer_0[2170] = in[213]; 
    assign layer_0[2171] = ~(in[67] ^ in[165]); 
    assign layer_0[2172] = ~(in[58] ^ in[70]); 
    assign layer_0[2173] = in[197]; 
    assign layer_0[2174] = ~(in[140] | in[156]); 
    assign layer_0[2175] = in[86] & ~in[25]; 
    assign layer_0[2176] = ~(in[5] | in[6]); 
    assign layer_0[2177] = ~in[150] | (in[92] & in[150]); 
    assign layer_0[2178] = in[215] & ~in[45]; 
    assign layer_0[2179] = ~(in[27] | in[191]); 
    assign layer_0[2180] = ~(in[89] ^ in[75]); 
    assign layer_0[2181] = in[119] ^ in[133]; 
    assign layer_0[2182] = in[115]; 
    assign layer_0[2183] = ~(in[6] | in[193]); 
    assign layer_0[2184] = 1'b1; 
    assign layer_0[2185] = ~in[178]; 
    assign layer_0[2186] = in[143] | in[194]; 
    assign layer_0[2187] = in[178]; 
    assign layer_0[2188] = in[56]; 
    assign layer_0[2189] = ~(in[185] ^ in[230]); 
    assign layer_0[2190] = ~(in[251] | in[22]); 
    assign layer_0[2191] = ~(in[90] ^ in[108]); 
    assign layer_0[2192] = ~(in[95] ^ in[5]); 
    assign layer_0[2193] = ~(in[183] & in[59]); 
    assign layer_0[2194] = ~(in[97] | in[249]); 
    assign layer_0[2195] = in[103] ^ in[134]; 
    assign layer_0[2196] = in[153] ^ in[123]; 
    assign layer_0[2197] = ~(in[22] ^ in[226]); 
    assign layer_0[2198] = ~in[29]; 
    assign layer_0[2199] = in[233] ^ in[78]; 
    assign layer_0[2200] = ~(in[100] | in[114]); 
    assign layer_0[2201] = ~in[140]; 
    assign layer_0[2202] = in[19] & ~in[146]; 
    assign layer_0[2203] = in[234] ^ in[196]; 
    assign layer_0[2204] = in[219] ^ in[73]; 
    assign layer_0[2205] = ~in[72] | (in[10] & in[72]); 
    assign layer_0[2206] = ~(in[109] ^ in[115]); 
    assign layer_0[2207] = in[170] & ~in[247]; 
    assign layer_0[2208] = in[133] & ~in[22]; 
    assign layer_0[2209] = in[148] | in[166]; 
    assign layer_0[2210] = ~(in[219] ^ in[123]); 
    assign layer_0[2211] = ~(in[50] ^ in[78]); 
    assign layer_0[2212] = in[87] & ~in[92]; 
    assign layer_0[2213] = ~(in[198] | in[5]); 
    assign layer_0[2214] = in[157] | in[143]; 
    assign layer_0[2215] = ~in[100] | (in[100] & in[157]); 
    assign layer_0[2216] = ~(in[143] | in[6]); 
    assign layer_0[2217] = in[216] & ~in[251]; 
    assign layer_0[2218] = in[137]; 
    assign layer_0[2219] = ~(in[76] ^ in[78]); 
    assign layer_0[2220] = in[90] | in[83]; 
    assign layer_0[2221] = ~(in[38] | in[242]); 
    assign layer_0[2222] = ~(in[56] ^ in[94]); 
    assign layer_0[2223] = ~in[147]; 
    assign layer_0[2224] = ~(in[97] & in[121]); 
    assign layer_0[2225] = in[165] ^ in[163]; 
    assign layer_0[2226] = ~(in[122] ^ in[138]); 
    assign layer_0[2227] = ~(in[74] ^ in[43]); 
    assign layer_0[2228] = in[200] ^ in[167]; 
    assign layer_0[2229] = in[181] ^ in[217]; 
    assign layer_0[2230] = ~(in[132] ^ in[149]); 
    assign layer_0[2231] = in[93] ^ in[91]; 
    assign layer_0[2232] = ~(in[197] | in[198]); 
    assign layer_0[2233] = in[89] ^ in[59]; 
    assign layer_0[2234] = in[167]; 
    assign layer_0[2235] = ~in[109] | (in[109] & in[232]); 
    assign layer_0[2236] = ~(in[87] ^ in[40]); 
    assign layer_0[2237] = ~in[132] | (in[11] & in[132]); 
    assign layer_0[2238] = in[62] ^ in[30]; 
    assign layer_0[2239] = ~(in[39] | in[55]); 
    assign layer_0[2240] = ~(in[130] | in[148]); 
    assign layer_0[2241] = ~in[130] | (in[170] & in[130]); 
    assign layer_0[2242] = ~(in[246] | in[215]); 
    assign layer_0[2243] = in[154] | in[99]; 
    assign layer_0[2244] = ~(in[57] ^ in[103]); 
    assign layer_0[2245] = ~in[250] | (in[250] & in[74]); 
    assign layer_0[2246] = ~(in[5] ^ in[139]); 
    assign layer_0[2247] = in[182] & ~in[170]; 
    assign layer_0[2248] = in[104] & ~in[109]; 
    assign layer_0[2249] = in[149] | in[236]; 
    assign layer_0[2250] = in[143] | in[73]; 
    assign layer_0[2251] = ~(in[167] | in[165]); 
    assign layer_0[2252] = in[170] & ~in[112]; 
    assign layer_0[2253] = ~(in[57] | in[25]); 
    assign layer_0[2254] = in[92] ^ in[94]; 
    assign layer_0[2255] = in[121] ^ in[22]; 
    assign layer_0[2256] = ~in[246] | (in[214] & in[246]); 
    assign layer_0[2257] = ~(in[26] | in[52]); 
    assign layer_0[2258] = ~in[142]; 
    assign layer_0[2259] = ~(in[35] | in[188]); 
    assign layer_0[2260] = ~in[231] | (in[231] & in[105]); 
    assign layer_0[2261] = ~(in[110] | in[137]); 
    assign layer_0[2262] = ~in[9]; 
    assign layer_0[2263] = in[152] ^ in[121]; 
    assign layer_0[2264] = in[119] ^ in[154]; 
    assign layer_0[2265] = ~(in[77] ^ in[44]); 
    assign layer_0[2266] = in[26] ^ in[209]; 
    assign layer_0[2267] = ~(in[107] ^ in[139]); 
    assign layer_0[2268] = ~in[124]; 
    assign layer_0[2269] = in[6]; 
    assign layer_0[2270] = in[46] ^ in[92]; 
    assign layer_0[2271] = ~in[102] | (in[102] & in[104]); 
    assign layer_0[2272] = in[74] ^ in[77]; 
    assign layer_0[2273] = ~(in[88] & in[183]); 
    assign layer_0[2274] = in[208] | in[5]; 
    assign layer_0[2275] = ~(in[146] ^ in[66]); 
    assign layer_0[2276] = ~(in[140] | in[49]); 
    assign layer_0[2277] = in[98] | in[180]; 
    assign layer_0[2278] = ~in[102] | (in[102] & in[90]); 
    assign layer_0[2279] = in[105] ^ in[183]; 
    assign layer_0[2280] = in[166] & ~in[245]; 
    assign layer_0[2281] = ~(in[100] | in[42]); 
    assign layer_0[2282] = ~in[135] | (in[135] & in[141]); 
    assign layer_0[2283] = in[194] ^ in[44]; 
    assign layer_0[2284] = ~(in[138] | in[23]); 
    assign layer_0[2285] = ~(in[47] | in[143]); 
    assign layer_0[2286] = ~in[134] | (in[131] & in[134]); 
    assign layer_0[2287] = in[168] & ~in[130]; 
    assign layer_0[2288] = ~(in[106] | in[219]); 
    assign layer_0[2289] = in[212] | in[135]; 
    assign layer_0[2290] = ~(in[146] ^ in[164]); 
    assign layer_0[2291] = in[188] & ~in[38]; 
    assign layer_0[2292] = ~(in[163] | in[177]); 
    assign layer_0[2293] = in[137] & ~in[139]; 
    assign layer_0[2294] = ~in[126]; 
    assign layer_0[2295] = in[244] ^ in[247]; 
    assign layer_0[2296] = in[39] ^ in[201]; 
    assign layer_0[2297] = in[155] | in[170]; 
    assign layer_0[2298] = in[82] | in[148]; 
    assign layer_0[2299] = in[248] | in[166]; 
    assign layer_0[2300] = ~(in[135] ^ in[166]); 
    assign layer_0[2301] = ~(in[101] ^ in[114]); 
    assign layer_0[2302] = ~in[117]; 
    assign layer_0[2303] = in[41] ^ in[171]; 
    assign layer_0[2304] = ~(in[112] | in[241]); 
    assign layer_0[2305] = in[63] | in[130]; 
    assign layer_0[2306] = in[168] & ~in[40]; 
    assign layer_0[2307] = ~(in[185] ^ in[37]); 
    assign layer_0[2308] = in[76] ^ in[72]; 
    assign layer_0[2309] = in[156] ^ in[203]; 
    assign layer_0[2310] = ~in[245] | (in[245] & in[196]); 
    assign layer_0[2311] = in[57]; 
    assign layer_0[2312] = in[185] & ~in[215]; 
    assign layer_0[2313] = in[7] ^ in[197]; 
    assign layer_0[2314] = ~in[34]; 
    assign layer_0[2315] = ~(in[129] ^ in[115]); 
    assign layer_0[2316] = ~(in[108] | in[125]); 
    assign layer_0[2317] = in[165] | in[146]; 
    assign layer_0[2318] = in[181] ^ in[99]; 
    assign layer_0[2319] = ~in[58] | (in[58] & in[218]); 
    assign layer_0[2320] = ~(in[42] ^ in[89]); 
    assign layer_0[2321] = ~(in[36] ^ in[195]); 
    assign layer_0[2322] = in[70] ^ in[83]; 
    assign layer_0[2323] = ~in[168] | (in[229] & in[168]); 
    assign layer_0[2324] = ~in[78]; 
    assign layer_0[2325] = in[9] ^ in[221]; 
    assign layer_0[2326] = in[139] & in[153]; 
    assign layer_0[2327] = in[163]; 
    assign layer_0[2328] = in[199]; 
    assign layer_0[2329] = in[178] | in[34]; 
    assign layer_0[2330] = in[98] | in[110]; 
    assign layer_0[2331] = ~in[83] | (in[83] & in[97]); 
    assign layer_0[2332] = ~in[247] | (in[247] & in[135]); 
    assign layer_0[2333] = ~(in[113] ^ in[119]); 
    assign layer_0[2334] = ~(in[211] ^ in[76]); 
    assign layer_0[2335] = in[24] | in[192]; 
    assign layer_0[2336] = ~in[129] | (in[10] & in[129]); 
    assign layer_0[2337] = ~(in[123] ^ in[152]); 
    assign layer_0[2338] = in[221] ^ in[212]; 
    assign layer_0[2339] = in[184] ^ in[230]; 
    assign layer_0[2340] = ~(in[154] | in[93]); 
    assign layer_0[2341] = in[197] & ~in[150]; 
    assign layer_0[2342] = ~(in[25] | in[44]); 
    assign layer_0[2343] = ~(in[40] | in[56]); 
    assign layer_0[2344] = in[172] ^ in[74]; 
    assign layer_0[2345] = ~(in[156] | in[75]); 
    assign layer_0[2346] = in[120] ^ in[171]; 
    assign layer_0[2347] = ~(in[82] | in[210]); 
    assign layer_0[2348] = ~(in[132] | in[10]); 
    assign layer_0[2349] = ~(in[131] ^ in[117]); 
    assign layer_0[2350] = ~(in[134] ^ in[132]); 
    assign layer_0[2351] = in[199] ^ in[218]; 
    assign layer_0[2352] = in[156] & ~in[206]; 
    assign layer_0[2353] = ~(in[22] ^ in[108]); 
    assign layer_0[2354] = in[212] ^ in[245]; 
    assign layer_0[2355] = ~(in[236] & in[128]); 
    assign layer_0[2356] = in[202] ^ in[99]; 
    assign layer_0[2357] = in[69] ^ in[23]; 
    assign layer_0[2358] = ~(in[213] ^ in[228]); 
    assign layer_0[2359] = ~(in[244] | in[79]); 
    assign layer_0[2360] = ~in[118]; 
    assign layer_0[2361] = in[42] | in[39]; 
    assign layer_0[2362] = ~(in[227] ^ in[247]); 
    assign layer_0[2363] = in[97] & ~in[120]; 
    assign layer_0[2364] = in[179] ^ in[53]; 
    assign layer_0[2365] = ~in[212] | (in[212] & in[17]); 
    assign layer_0[2366] = ~in[152]; 
    assign layer_0[2367] = ~(in[165] ^ in[135]); 
    assign layer_0[2368] = in[103] ^ in[241]; 
    assign layer_0[2369] = ~(in[58] ^ in[11]); 
    assign layer_0[2370] = ~in[155] | (in[155] & in[196]); 
    assign layer_0[2371] = in[201] & in[219]; 
    assign layer_0[2372] = in[249] | in[220]; 
    assign layer_0[2373] = ~in[9]; 
    assign layer_0[2374] = in[215]; 
    assign layer_0[2375] = in[156] ^ in[138]; 
    assign layer_0[2376] = in[251] | in[190]; 
    assign layer_0[2377] = in[92] ^ in[90]; 
    assign layer_0[2378] = ~(in[73] ^ in[91]); 
    assign layer_0[2379] = in[51]; 
    assign layer_0[2380] = ~(in[173] | in[241]); 
    assign layer_0[2381] = ~(in[7] ^ in[69]); 
    assign layer_0[2382] = ~(in[106] | in[51]); 
    assign layer_0[2383] = in[118] | in[101]; 
    assign layer_0[2384] = ~in[25] | (in[25] & in[88]); 
    assign layer_0[2385] = in[125] ^ in[169]; 
    assign layer_0[2386] = in[104] ^ in[197]; 
    assign layer_0[2387] = ~(in[54] ^ in[99]); 
    assign layer_0[2388] = ~in[55] | (in[68] & in[55]); 
    assign layer_0[2389] = ~in[169] | (in[59] & in[169]); 
    assign layer_0[2390] = ~(in[108] ^ in[106]); 
    assign layer_0[2391] = ~in[27]; 
    assign layer_0[2392] = ~(in[106] | in[57]); 
    assign layer_0[2393] = ~(in[72] & in[191]); 
    assign layer_0[2394] = ~(in[203] ^ in[173]); 
    assign layer_0[2395] = in[220]; 
    assign layer_0[2396] = ~(in[22] ^ in[214]); 
    assign layer_0[2397] = in[153] & ~in[196]; 
    assign layer_0[2398] = in[242] ^ in[66]; 
    assign layer_0[2399] = ~in[167] | (in[77] & in[167]); 
    assign layer_0[2400] = in[90]; 
    assign layer_0[2401] = in[72] & ~in[11]; 
    assign layer_0[2402] = ~(in[40] ^ in[113]); 
    assign layer_0[2403] = in[249]; 
    assign layer_0[2404] = ~in[58] | (in[58] & in[85]); 
    assign layer_0[2405] = in[104] | in[118]; 
    assign layer_0[2406] = in[118]; 
    assign layer_0[2407] = in[61] ^ in[92]; 
    assign layer_0[2408] = in[153] ^ in[118]; 
    assign layer_0[2409] = in[194] | in[219]; 
    assign layer_0[2410] = in[154]; 
    assign layer_0[2411] = in[39] & ~in[219]; 
    assign layer_0[2412] = in[106] ^ in[163]; 
    assign layer_0[2413] = in[101]; 
    assign layer_0[2414] = in[232] & ~in[10]; 
    assign layer_0[2415] = in[231] ^ in[200]; 
    assign layer_0[2416] = ~(in[94] ^ in[50]); 
    assign layer_0[2417] = ~in[110]; 
    assign layer_0[2418] = ~in[235]; 
    assign layer_0[2419] = ~(in[123] | in[140]); 
    assign layer_0[2420] = in[148]; 
    assign layer_0[2421] = ~(in[149] ^ in[147]); 
    assign layer_0[2422] = in[214]; 
    assign layer_0[2423] = ~(in[169] ^ in[149]); 
    assign layer_0[2424] = ~(in[78] ^ in[21]); 
    assign layer_0[2425] = in[226] ^ in[245]; 
    assign layer_0[2426] = ~(in[37] ^ in[73]); 
    assign layer_0[2427] = in[58] ^ in[111]; 
    assign layer_0[2428] = ~in[187]; 
    assign layer_0[2429] = in[120]; 
    assign layer_0[2430] = ~(in[189] | in[251]); 
    assign layer_0[2431] = in[234]; 
    assign layer_0[2432] = in[139] | in[106]; 
    assign layer_0[2433] = ~(in[170] ^ in[233]); 
    assign layer_0[2434] = ~(in[148] ^ in[180]); 
    assign layer_0[2435] = in[251] ^ in[204]; 
    assign layer_0[2436] = ~(in[165] | in[163]); 
    assign layer_0[2437] = ~in[133] | (in[133] & in[74]); 
    assign layer_0[2438] = in[44]; 
    assign layer_0[2439] = ~in[201] | (in[201] & in[55]); 
    assign layer_0[2440] = ~in[137] | (in[187] & in[137]); 
    assign layer_0[2441] = in[120] ^ in[74]; 
    assign layer_0[2442] = in[116] ^ in[129]; 
    assign layer_0[2443] = in[93] ^ in[91]; 
    assign layer_0[2444] = in[22] ^ in[36]; 
    assign layer_0[2445] = ~(in[73] ^ in[77]); 
    assign layer_0[2446] = in[54] & in[86]; 
    assign layer_0[2447] = ~(in[21] ^ in[143]); 
    assign layer_0[2448] = ~in[132]; 
    assign layer_0[2449] = in[237] & ~in[204]; 
    assign layer_0[2450] = ~(in[132] ^ in[146]); 
    assign layer_0[2451] = in[195] ^ in[187]; 
    assign layer_0[2452] = in[133]; 
    assign layer_0[2453] = in[211]; 
    assign layer_0[2454] = ~(in[166] | in[131]); 
    assign layer_0[2455] = in[90] | in[45]; 
    assign layer_0[2456] = ~(in[189] & in[222]); 
    assign layer_0[2457] = ~(in[114] ^ in[186]); 
    assign layer_0[2458] = in[38] ^ in[195]; 
    assign layer_0[2459] = in[217] & ~in[107]; 
    assign layer_0[2460] = ~in[154] | (in[212] & in[154]); 
    assign layer_0[2461] = ~(in[107] ^ in[89]); 
    assign layer_0[2462] = ~in[248]; 
    assign layer_0[2463] = in[29] & ~in[114]; 
    assign layer_0[2464] = ~(in[69] ^ in[89]); 
    assign layer_0[2465] = ~(in[122] ^ in[74]); 
    assign layer_0[2466] = ~(in[100] ^ in[86]); 
    assign layer_0[2467] = in[131] | in[148]; 
    assign layer_0[2468] = in[67] ^ in[87]; 
    assign layer_0[2469] = in[28] ^ in[8]; 
    assign layer_0[2470] = ~in[247]; 
    assign layer_0[2471] = in[250] ^ in[248]; 
    assign layer_0[2472] = ~(in[143] ^ in[196]); 
    assign layer_0[2473] = ~(in[145] ^ in[147]); 
    assign layer_0[2474] = in[249] & ~in[159]; 
    assign layer_0[2475] = ~(in[133] | in[162]); 
    assign layer_0[2476] = in[71] ^ in[85]; 
    assign layer_0[2477] = in[108] & ~in[79]; 
    assign layer_0[2478] = ~(in[101] ^ in[70]); 
    assign layer_0[2479] = in[26] & ~in[72]; 
    assign layer_0[2480] = in[212] ^ in[227]; 
    assign layer_0[2481] = ~(in[142] | in[11]); 
    assign layer_0[2482] = in[155] & ~in[27]; 
    assign layer_0[2483] = in[184] | in[212]; 
    assign layer_0[2484] = in[164] & ~in[12]; 
    assign layer_0[2485] = ~(in[73] ^ in[42]); 
    assign layer_0[2486] = in[118] ^ in[90]; 
    assign layer_0[2487] = ~(in[109] ^ in[91]); 
    assign layer_0[2488] = ~(in[172] | in[126]); 
    assign layer_0[2489] = in[168] & ~in[203]; 
    assign layer_0[2490] = in[219] ^ in[189]; 
    assign layer_0[2491] = ~(in[136] ^ in[187]); 
    assign layer_0[2492] = ~(in[163] ^ in[181]); 
    assign layer_0[2493] = ~(in[180] ^ in[215]); 
    assign layer_0[2494] = ~in[81]; 
    assign layer_0[2495] = ~(in[68] | in[68]); 
    assign layer_0[2496] = ~(in[24] ^ in[71]); 
    assign layer_0[2497] = ~(in[79] | in[218]); 
    assign layer_0[2498] = ~in[153] | (in[180] & in[153]); 
    assign layer_0[2499] = ~(in[178] ^ in[196]); 
    assign layer_0[2500] = in[242]; 
    assign layer_0[2501] = ~(in[168] ^ in[251]); 
    assign layer_0[2502] = in[113] | in[114]; 
    assign layer_0[2503] = ~in[216] | (in[216] & in[244]); 
    assign layer_0[2504] = ~(in[53] ^ in[5]); 
    assign layer_0[2505] = ~in[119]; 
    assign layer_0[2506] = in[169] & ~in[196]; 
    assign layer_0[2507] = ~(in[215] | in[213]); 
    assign layer_0[2508] = ~(in[148] ^ in[165]); 
    assign layer_0[2509] = ~(in[53] | in[42]); 
    assign layer_0[2510] = ~in[153] | (in[153] & in[83]); 
    assign layer_0[2511] = ~in[103] | (in[134] & in[103]); 
    assign layer_0[2512] = ~(in[233] ^ in[165]); 
    assign layer_0[2513] = ~(in[85] ^ in[87]); 
    assign layer_0[2514] = ~(in[205] | in[195]); 
    assign layer_0[2515] = ~(in[77] | in[229]); 
    assign layer_0[2516] = ~(in[20] ^ in[235]); 
    assign layer_0[2517] = ~in[73] | (in[182] & in[73]); 
    assign layer_0[2518] = in[163] | in[146]; 
    assign layer_0[2519] = in[219] & ~in[114]; 
    assign layer_0[2520] = ~(in[173] & in[71]); 
    assign layer_0[2521] = ~(in[78] | in[108]); 
    assign layer_0[2522] = ~(in[11] ^ in[111]); 
    assign layer_0[2523] = ~in[220]; 
    assign layer_0[2524] = in[19] | in[141]; 
    assign layer_0[2525] = ~(in[139] ^ in[186]); 
    assign layer_0[2526] = ~in[132] | (in[130] & in[132]); 
    assign layer_0[2527] = in[60] | in[34]; 
    assign layer_0[2528] = ~(in[99] ^ in[167]); 
    assign layer_0[2529] = ~in[90]; 
    assign layer_0[2530] = ~in[147] | (in[147] & in[138]); 
    assign layer_0[2531] = in[228] ^ in[177]; 
    assign layer_0[2532] = in[196] & ~in[227]; 
    assign layer_0[2533] = in[119] & ~in[124]; 
    assign layer_0[2534] = ~(in[203] ^ in[248]); 
    assign layer_0[2535] = ~in[196] | (in[196] & in[12]); 
    assign layer_0[2536] = ~in[21]; 
    assign layer_0[2537] = in[106] ^ in[75]; 
    assign layer_0[2538] = in[24] | in[26]; 
    assign layer_0[2539] = in[30] | in[101]; 
    assign layer_0[2540] = ~(in[78] | in[228]); 
    assign layer_0[2541] = in[211] ^ in[196]; 
    assign layer_0[2542] = in[97] ^ in[99]; 
    assign layer_0[2543] = ~(in[139] | in[185]); 
    assign layer_0[2544] = ~(in[89] ^ in[138]); 
    assign layer_0[2545] = in[125] & ~in[148]; 
    assign layer_0[2546] = in[166] ^ in[120]; 
    assign layer_0[2547] = ~(in[232] ^ in[10]); 
    assign layer_0[2548] = in[136] ^ in[104]; 
    assign layer_0[2549] = in[100] ^ in[102]; 
    assign layer_0[2550] = in[38] ^ in[70]; 
    assign layer_0[2551] = ~(in[118] | in[25]); 
    assign layer_0[2552] = in[182] & ~in[76]; 
    assign layer_0[2553] = ~in[121] | (in[50] & in[121]); 
    assign layer_0[2554] = in[109] ^ in[170]; 
    assign layer_0[2555] = in[36]; 
    assign layer_0[2556] = in[189] ^ in[108]; 
    assign layer_0[2557] = in[99] ^ in[68]; 
    assign layer_0[2558] = in[143] & ~in[114]; 
    assign layer_0[2559] = ~(in[121] ^ in[123]); 
    // Layer 1 ============================================================
    assign out[0] = layer_0[56]; 
    assign out[1] = layer_0[258] ^ layer_0[1272]; 
    assign out[2] = layer_0[266]; 
    assign out[3] = ~(layer_0[1651] & layer_0[954]); 
    assign out[4] = ~layer_0[2264]; 
    assign out[5] = ~layer_0[1625]; 
    assign out[6] = ~(layer_0[512] & layer_0[358]); 
    assign out[7] = ~(layer_0[1461] | layer_0[2093]); 
    assign out[8] = layer_0[1187]; 
    assign out[9] = layer_0[1690]; 
    assign out[10] = layer_0[1641] ^ layer_0[1357]; 
    assign out[11] = ~(layer_0[751] ^ layer_0[1085]); 
    assign out[12] = ~(layer_0[1365] | layer_0[860]); 
    assign out[13] = ~layer_0[1574]; 
    assign out[14] = layer_0[1212]; 
    assign out[15] = ~layer_0[1274] | (layer_0[1274] & layer_0[792]); 
    assign out[16] = ~layer_0[322] | (layer_0[657] & layer_0[322]); 
    assign out[17] = ~(layer_0[2340] ^ layer_0[2551]); 
    assign out[18] = layer_0[1273] ^ layer_0[1724]; 
    assign out[19] = ~(layer_0[390] ^ layer_0[2526]); 
    assign out[20] = layer_0[969] & ~layer_0[1095]; 
    assign out[21] = ~layer_0[2263]; 
    assign out[22] = ~(layer_0[1281] ^ layer_0[982]); 
    assign out[23] = layer_0[924]; 
    assign out[24] = layer_0[709] & layer_0[2123]; 
    assign out[25] = ~layer_0[555] | (layer_0[555] & layer_0[217]); 
    assign out[26] = layer_0[268] ^ layer_0[2234]; 
    assign out[27] = ~layer_0[2357]; 
    assign out[28] = layer_0[619] & layer_0[2498]; 
    assign out[29] = ~layer_0[769]; 
    assign out[30] = ~layer_0[1412] | (layer_0[216] & layer_0[1412]); 
    assign out[31] = ~layer_0[2372]; 
    assign out[32] = layer_0[1883] & ~layer_0[1488]; 
    assign out[33] = layer_0[2292] ^ layer_0[2053]; 
    assign out[34] = ~(layer_0[814] | layer_0[2403]); 
    assign out[35] = layer_0[1619]; 
    assign out[36] = layer_0[222]; 
    assign out[37] = layer_0[2474] ^ layer_0[912]; 
    assign out[38] = layer_0[474] & ~layer_0[548]; 
    assign out[39] = ~layer_0[450] | (layer_0[1837] & layer_0[450]); 
    assign out[40] = layer_0[2241] ^ layer_0[2350]; 
    assign out[41] = ~(layer_0[29] ^ layer_0[870]); 
    assign out[42] = layer_0[740] & ~layer_0[2033]; 
    assign out[43] = layer_0[660]; 
    assign out[44] = layer_0[2260] ^ layer_0[16]; 
    assign out[45] = layer_0[687] ^ layer_0[187]; 
    assign out[46] = ~layer_0[309]; 
    assign out[47] = ~layer_0[1594]; 
    assign out[48] = layer_0[1063] & ~layer_0[585]; 
    assign out[49] = ~(layer_0[2095] ^ layer_0[786]); 
    assign out[50] = ~layer_0[1672]; 
    assign out[51] = layer_0[935] & ~layer_0[1176]; 
    assign out[52] = layer_0[2544]; 
    assign out[53] = ~(layer_0[1530] | layer_0[861]); 
    assign out[54] = layer_0[1242] & layer_0[461]; 
    assign out[55] = layer_0[1445] | layer_0[1808]; 
    assign out[56] = layer_0[559] ^ layer_0[1009]; 
    assign out[57] = ~layer_0[267]; 
    assign out[58] = layer_0[365] ^ layer_0[1498]; 
    assign out[59] = layer_0[903] & ~layer_0[2255]; 
    assign out[60] = ~(layer_0[2078] | layer_0[1802]); 
    assign out[61] = layer_0[271] & layer_0[215]; 
    assign out[62] = layer_0[794] & layer_0[770]; 
    assign out[63] = ~(layer_0[856] ^ layer_0[303]); 
    assign out[64] = ~layer_0[1809]; 
    assign out[65] = ~(layer_0[41] | layer_0[1796]); 
    assign out[66] = ~(layer_0[59] ^ layer_0[568]); 
    assign out[67] = ~layer_0[869]; 
    assign out[68] = ~(layer_0[398] ^ layer_0[2279]); 
    assign out[69] = layer_0[468] & ~layer_0[1145]; 
    assign out[70] = ~layer_0[531]; 
    assign out[71] = layer_0[524] ^ layer_0[836]; 
    assign out[72] = ~layer_0[1158]; 
    assign out[73] = layer_0[2167]; 
    assign out[74] = ~(layer_0[1065] ^ layer_0[1236]); 
    assign out[75] = layer_0[1591] ^ layer_0[272]; 
    assign out[76] = layer_0[48]; 
    assign out[77] = layer_0[621] ^ layer_0[1277]; 
    assign out[78] = ~(layer_0[948] & layer_0[1379]); 
    assign out[79] = ~(layer_0[50] | layer_0[1806]); 
    assign out[80] = layer_0[1951]; 
    assign out[81] = layer_0[2516] & layer_0[1586]; 
    assign out[82] = ~(layer_0[2287] | layer_0[577]); 
    assign out[83] = ~(layer_0[102] ^ layer_0[1303]); 
    assign out[84] = layer_0[1109] ^ layer_0[2185]; 
    assign out[85] = ~layer_0[1867]; 
    assign out[86] = ~(layer_0[12] ^ layer_0[2031]); 
    assign out[87] = layer_0[1816] & ~layer_0[435]; 
    assign out[88] = ~(layer_0[1841] ^ layer_0[183]); 
    assign out[89] = ~layer_0[2195]; 
    assign out[90] = layer_0[313] & ~layer_0[487]; 
    assign out[91] = ~(layer_0[1447] & layer_0[1030]); 
    assign out[92] = layer_0[991] ^ layer_0[575]; 
    assign out[93] = layer_0[1994] ^ layer_0[1992]; 
    assign out[94] = ~(layer_0[1258] & layer_0[1991]); 
    assign out[95] = ~(layer_0[1914] ^ layer_0[1123]); 
    assign out[96] = layer_0[2226] & ~layer_0[806]; 
    assign out[97] = ~(layer_0[1204] ^ layer_0[2477]); 
    assign out[98] = layer_0[1356]; 
    assign out[99] = ~(layer_0[578] ^ layer_0[227]); 
    assign out[100] = layer_0[1430] ^ layer_0[1861]; 
    assign out[101] = ~layer_0[1108] | (layer_0[5] & layer_0[1108]); 
    assign out[102] = layer_0[386] & layer_0[2518]; 
    assign out[103] = layer_0[929] & layer_0[1814]; 
    assign out[104] = ~(layer_0[444] ^ layer_0[1372]); 
    assign out[105] = layer_0[66]; 
    assign out[106] = layer_0[2467] & layer_0[1917]; 
    assign out[107] = layer_0[1294] ^ layer_0[388]; 
    assign out[108] = ~layer_0[1970] | (layer_0[2055] & layer_0[1970]); 
    assign out[109] = layer_0[2131] & ~layer_0[644]; 
    assign out[110] = layer_0[2013]; 
    assign out[111] = ~layer_0[2074]; 
    assign out[112] = ~(layer_0[2331] ^ layer_0[1064]); 
    assign out[113] = ~layer_0[1453] | (layer_0[1453] & layer_0[391]); 
    assign out[114] = layer_0[1790] & ~layer_0[329]; 
    assign out[115] = ~layer_0[1956]; 
    assign out[116] = layer_0[2134] ^ layer_0[2361]; 
    assign out[117] = layer_0[1972] | layer_0[1930]; 
    assign out[118] = layer_0[400] & layer_0[682]; 
    assign out[119] = ~(layer_0[781] ^ layer_0[181]); 
    assign out[120] = ~layer_0[1953] | (layer_0[2047] & layer_0[1953]); 
    assign out[121] = layer_0[810]; 
    assign out[122] = layer_0[2157] | layer_0[1450]; 
    assign out[123] = ~layer_0[679] | (layer_0[368] & layer_0[679]); 
    assign out[124] = layer_0[2105]; 
    assign out[125] = ~layer_0[1546] | (layer_0[1546] & layer_0[1124]); 
    assign out[126] = ~layer_0[1614]; 
    assign out[127] = layer_0[2066] ^ layer_0[2464]; 
    assign out[128] = layer_0[1691]; 
    assign out[129] = layer_0[764] | layer_0[1940]; 
    assign out[130] = ~(layer_0[1709] ^ layer_0[85]); 
    assign out[131] = ~(layer_0[1196] | layer_0[1974]); 
    assign out[132] = ~(layer_0[1610] | layer_0[2005]); 
    assign out[133] = layer_0[1333]; 
    assign out[134] = layer_0[2229]; 
    assign out[135] = ~(layer_0[2112] ^ layer_0[2048]); 
    assign out[136] = layer_0[1103] ^ layer_0[2107]; 
    assign out[137] = ~layer_0[22]; 
    assign out[138] = layer_0[456] ^ layer_0[2555]; 
    assign out[139] = layer_0[295]; 
    assign out[140] = layer_0[2307]; 
    assign out[141] = ~(layer_0[1257] ^ layer_0[1159]); 
    assign out[142] = layer_0[276] ^ layer_0[2189]; 
    assign out[143] = ~(layer_0[1471] ^ layer_0[1249]); 
    assign out[144] = layer_0[2197] & ~layer_0[1229]; 
    assign out[145] = layer_0[1409] | layer_0[983]; 
    assign out[146] = ~(layer_0[721] ^ layer_0[202]); 
    assign out[147] = ~(layer_0[1153] | layer_0[418]); 
    assign out[148] = layer_0[35] | layer_0[988]; 
    assign out[149] = ~layer_0[787] | (layer_0[123] & layer_0[787]); 
    assign out[150] = layer_0[1731] & ~layer_0[485]; 
    assign out[151] = layer_0[164] ^ layer_0[2086]; 
    assign out[152] = ~layer_0[2084]; 
    assign out[153] = ~layer_0[1937]; 
    assign out[154] = layer_0[2158] & ~layer_0[415]; 
    assign out[155] = layer_0[111]; 
    assign out[156] = layer_0[973] ^ layer_0[622]; 
    assign out[157] = ~(layer_0[2288] ^ layer_0[2510]); 
    assign out[158] = ~(layer_0[2284] ^ layer_0[1435]); 
    assign out[159] = layer_0[1702] & layer_0[976]; 
    assign out[160] = ~(layer_0[1053] ^ layer_0[1636]); 
    assign out[161] = ~layer_0[638] | (layer_0[1033] & layer_0[638]); 
    assign out[162] = layer_0[2504] & ~layer_0[327]; 
    assign out[163] = layer_0[2483] & ~layer_0[737]; 
    assign out[164] = ~layer_0[1380]; 
    assign out[165] = ~layer_0[1089] | (layer_0[1089] & layer_0[1205]); 
    assign out[166] = layer_0[167] & layer_0[1499]; 
    assign out[167] = layer_0[325] & ~layer_0[1888]; 
    assign out[168] = ~(layer_0[586] & layer_0[1282]); 
    assign out[169] = ~layer_0[2493]; 
    assign out[170] = layer_0[2015]; 
    assign out[171] = ~(layer_0[2293] ^ layer_0[1349]); 
    assign out[172] = ~(layer_0[1767] ^ layer_0[1587]); 
    assign out[173] = ~layer_0[616]; 
    assign out[174] = ~(layer_0[1759] ^ layer_0[2538]); 
    assign out[175] = ~(layer_0[1364] ^ layer_0[2079]); 
    assign out[176] = ~(layer_0[767] ^ layer_0[196]); 
    assign out[177] = layer_0[1517] & layer_0[1567]; 
    assign out[178] = layer_0[126] ^ layer_0[2369]; 
    assign out[179] = ~(layer_0[985] & layer_0[2057]); 
    assign out[180] = layer_0[1935] ^ layer_0[1174]; 
    assign out[181] = layer_0[752]; 
    assign out[182] = layer_0[475] ^ layer_0[551]; 
    assign out[183] = ~(layer_0[2318] | layer_0[374]); 
    assign out[184] = ~layer_0[1375] | (layer_0[1851] & layer_0[1375]); 
    assign out[185] = ~(layer_0[2114] ^ layer_0[2299]); 
    assign out[186] = ~layer_0[446]; 
    assign out[187] = ~layer_0[1723] | (layer_0[1316] & layer_0[1723]); 
    assign out[188] = layer_0[1125] | layer_0[38]; 
    assign out[189] = ~(layer_0[945] ^ layer_0[1162]); 
    assign out[190] = layer_0[1348] ^ layer_0[1857]; 
    assign out[191] = layer_0[1466] & ~layer_0[1134]; 
    assign out[192] = layer_0[1798] & layer_0[1317]; 
    assign out[193] = layer_0[2465] & layer_0[1620]; 
    assign out[194] = layer_0[2458] ^ layer_0[1795]; 
    assign out[195] = layer_0[2002] & layer_0[1363]; 
    assign out[196] = layer_0[344]; 
    assign out[197] = ~(layer_0[766] | layer_0[727]); 
    assign out[198] = layer_0[1458] | layer_0[2371]; 
    assign out[199] = ~(layer_0[1697] | layer_0[1289]); 
    assign out[200] = layer_0[292]; 
    assign out[201] = ~layer_0[529] | (layer_0[105] & layer_0[529]); 
    assign out[202] = ~(layer_0[1407] ^ layer_0[1561]); 
    assign out[203] = layer_0[1338] & layer_0[1276]; 
    assign out[204] = layer_0[2382] ^ layer_0[1329]; 
    assign out[205] = ~layer_0[2534]; 
    assign out[206] = layer_0[2421] & layer_0[55]; 
    assign out[207] = layer_0[2281] & layer_0[262]; 
    assign out[208] = layer_0[1853] & layer_0[488]; 
    assign out[209] = ~(layer_0[1077] | layer_0[937]); 
    assign out[210] = ~layer_0[824]; 
    assign out[211] = ~layer_0[67] | (layer_0[67] & layer_0[1668]); 
    assign out[212] = layer_0[265] & ~layer_0[649]; 
    assign out[213] = ~layer_0[2423]; 
    assign out[214] = layer_0[1746] & ~layer_0[838]; 
    assign out[215] = layer_0[205]; 
    assign out[216] = layer_0[1783] ^ layer_0[1496]; 
    assign out[217] = ~(layer_0[1040] ^ layer_0[382]); 
    assign out[218] = layer_0[1484] ^ layer_0[1128]; 
    assign out[219] = layer_0[60] & ~layer_0[748]; 
    assign out[220] = layer_0[1474]; 
    assign out[221] = layer_0[1200] & ~layer_0[330]; 
    assign out[222] = ~(layer_0[1577] | layer_0[2072]); 
    assign out[223] = layer_0[2408] & ~layer_0[1221]; 
    assign out[224] = layer_0[1490] & layer_0[1015]; 
    assign out[225] = ~(layer_0[286] ^ layer_0[19]); 
    assign out[226] = ~(layer_0[1737] ^ layer_0[1889]); 
    assign out[227] = layer_0[1102] ^ layer_0[1933]; 
    assign out[228] = layer_0[778] & layer_0[518]; 
    assign out[229] = layer_0[2006] ^ layer_0[2321]; 
    assign out[230] = layer_0[651] ^ layer_0[1791]; 
    assign out[231] = layer_0[2426] ^ layer_0[350]; 
    assign out[232] = layer_0[839]; 
    assign out[233] = layer_0[2308] & ~layer_0[404]; 
    assign out[234] = layer_0[930] & layer_0[731]; 
    assign out[235] = ~layer_0[2270]; 
    assign out[236] = layer_0[1446] & ~layer_0[1824]; 
    assign out[237] = ~layer_0[826]; 
    assign out[238] = layer_0[1703] & ~layer_0[1870]; 
    assign out[239] = layer_0[706] | layer_0[1769]; 
    assign out[240] = ~(layer_0[225] | layer_0[332]); 
    assign out[241] = layer_0[746]; 
    assign out[242] = ~(layer_0[891] ^ layer_0[2553]); 
    assign out[243] = layer_0[1395] ^ layer_0[1149]; 
    assign out[244] = ~(layer_0[1394] ^ layer_0[1885]); 
    assign out[245] = layer_0[561] & layer_0[277]; 
    assign out[246] = ~(layer_0[1710] ^ layer_0[14]); 
    assign out[247] = ~layer_0[2243]; 
    assign out[248] = layer_0[2490]; 
    assign out[249] = ~layer_0[2172]; 
    assign out[250] = layer_0[2379] ^ layer_0[1195]; 
    assign out[251] = ~layer_0[335]; 
    assign out[252] = ~(layer_0[1084] ^ layer_0[219]); 
    assign out[253] = layer_0[2271] & ~layer_0[516]; 
    assign out[254] = ~(layer_0[441] ^ layer_0[845]); 
    assign out[255] = layer_0[2061] ^ layer_0[1314]; 
    assign out[256] = ~(layer_0[890] | layer_0[999]); 
    assign out[257] = layer_0[805]; 
    assign out[258] = layer_0[2155]; 
    assign out[259] = ~layer_0[2468] | (layer_0[2531] & layer_0[2468]); 
    assign out[260] = layer_0[1502] ^ layer_0[1382]; 
    assign out[261] = layer_0[2310] & ~layer_0[1643]; 
    assign out[262] = layer_0[1540] ^ layer_0[1214]; 
    assign out[263] = ~(layer_0[734] ^ layer_0[341]); 
    assign out[264] = ~(layer_0[1818] & layer_0[379]); 
    assign out[265] = ~layer_0[34] | (layer_0[1683] & layer_0[34]); 
    assign out[266] = layer_0[270] ^ layer_0[761]; 
    assign out[267] = layer_0[279] ^ layer_0[2054]; 
    assign out[268] = ~layer_0[2132] | (layer_0[2132] & layer_0[121]); 
    assign out[269] = ~layer_0[715]; 
    assign out[270] = layer_0[1341] ^ layer_0[2064]; 
    assign out[271] = ~(layer_0[245] & layer_0[784]); 
    assign out[272] = ~(layer_0[670] ^ layer_0[2007]); 
    assign out[273] = layer_0[1605] ^ layer_0[641]; 
    assign out[274] = layer_0[155] ^ layer_0[1649]; 
    assign out[275] = layer_0[1463] ^ layer_0[2135]; 
    assign out[276] = layer_0[96] ^ layer_0[627]; 
    assign out[277] = layer_0[1164] ^ layer_0[1927]; 
    assign out[278] = layer_0[1707] ^ layer_0[972]; 
    assign out[279] = layer_0[104] ^ layer_0[1126]; 
    assign out[280] = ~layer_0[1650]; 
    assign out[281] = layer_0[1830] ^ layer_0[895]; 
    assign out[282] = layer_0[81] & layer_0[264]; 
    assign out[283] = layer_0[1909] ^ layer_0[1464]; 
    assign out[284] = ~layer_0[351] | (layer_0[1460] & layer_0[351]); 
    assign out[285] = ~layer_0[1420]; 
    assign out[286] = layer_0[2368] ^ layer_0[1658]; 
    assign out[287] = layer_0[1952]; 
    assign out[288] = layer_0[17]; 
    assign out[289] = layer_0[931] ^ layer_0[1829]; 
    assign out[290] = layer_0[2303]; 
    assign out[291] = layer_0[355] ^ layer_0[1705]; 
    assign out[292] = ~(layer_0[694] | layer_0[1155]); 
    assign out[293] = layer_0[287] | layer_0[2558]; 
    assign out[294] = layer_0[1629]; 
    assign out[295] = ~(layer_0[635] ^ layer_0[1834]); 
    assign out[296] = layer_0[813] & ~layer_0[432]; 
    assign out[297] = layer_0[684]; 
    assign out[298] = layer_0[2339]; 
    assign out[299] = ~(layer_0[601] & layer_0[1414]); 
    assign out[300] = layer_0[148] ^ layer_0[1071]; 
    assign out[301] = layer_0[9] ^ layer_0[1288]; 
    assign out[302] = ~layer_0[2389] | (layer_0[2389] & layer_0[2479]); 
    assign out[303] = layer_0[1313] & ~layer_0[1189]; 
    assign out[304] = ~(layer_0[911] & layer_0[671]); 
    assign out[305] = ~(layer_0[28] ^ layer_0[1443]); 
    assign out[306] = layer_0[1508]; 
    assign out[307] = ~(layer_0[2449] ^ layer_0[1487]); 
    assign out[308] = ~(layer_0[686] ^ layer_0[850]); 
    assign out[309] = layer_0[2228]; 
    assign out[310] = layer_0[885] ^ layer_0[2384]; 
    assign out[311] = ~layer_0[2196]; 
    assign out[312] = ~(layer_0[724] ^ layer_0[1877]); 
    assign out[313] = ~(layer_0[274] ^ layer_0[708]); 
    assign out[314] = layer_0[2500] ^ layer_0[1104]; 
    assign out[315] = layer_0[2376] ^ layer_0[2395]; 
    assign out[316] = ~(layer_0[1262] ^ layer_0[1051]); 
    assign out[317] = layer_0[876] | layer_0[2147]; 
    assign out[318] = ~layer_0[174]; 
    assign out[319] = layer_0[395] & layer_0[1653]; 
    assign out[320] = layer_0[2166]; 
    assign out[321] = layer_0[1946] ^ layer_0[2001]; 
    assign out[322] = ~layer_0[793] | (layer_0[1986] & layer_0[793]); 
    assign out[323] = layer_0[943] | layer_0[51]; 
    assign out[324] = layer_0[1184] | layer_0[1961]; 
    assign out[325] = layer_0[1634] & layer_0[423]; 
    assign out[326] = ~layer_0[86] | (layer_0[1862] & layer_0[86]); 
    assign out[327] = ~(layer_0[502] ^ layer_0[128]); 
    assign out[328] = ~layer_0[1858] | (layer_0[232] & layer_0[1858]); 
    assign out[329] = layer_0[1451] | layer_0[2326]; 
    assign out[330] = ~(layer_0[816] & layer_0[558]); 
    assign out[331] = ~(layer_0[1058] ^ layer_0[293]); 
    assign out[332] = layer_0[1075]; 
    assign out[333] = ~layer_0[1425] | (layer_0[717] & layer_0[1425]); 
    assign out[334] = layer_0[371] | layer_0[950]; 
    assign out[335] = ~layer_0[926]; 
    assign out[336] = ~(layer_0[825] ^ layer_0[402]); 
    assign out[337] = ~layer_0[1810] | (layer_0[630] & layer_0[1810]); 
    assign out[338] = ~(layer_0[2163] ^ layer_0[302]); 
    assign out[339] = layer_0[2430] ^ layer_0[2523]; 
    assign out[340] = ~layer_0[1393]; 
    assign out[341] = ~layer_0[1863] | (layer_0[1863] & layer_0[1627]); 
    assign out[342] = ~(layer_0[243] ^ layer_0[2381]); 
    assign out[343] = ~layer_0[429]; 
    assign out[344] = layer_0[317] ^ layer_0[1993]; 
    assign out[345] = ~layer_0[2089]; 
    assign out[346] = ~(layer_0[981] & layer_0[743]); 
    assign out[347] = ~layer_0[2332] | (layer_0[1452] & layer_0[2332]); 
    assign out[348] = layer_0[757] ^ layer_0[1799]; 
    assign out[349] = layer_0[1304] ^ layer_0[1010]; 
    assign out[350] = ~(layer_0[854] ^ layer_0[1603]); 
    assign out[351] = layer_0[1390] ^ layer_0[1741]; 
    assign out[352] = layer_0[192]; 
    assign out[353] = layer_0[26] ^ layer_0[1589]; 
    assign out[354] = layer_0[1476] ^ layer_0[144]; 
    assign out[355] = ~(layer_0[2179] ^ layer_0[1081]); 
    assign out[356] = layer_0[1270] ^ layer_0[1087]; 
    assign out[357] = layer_0[2362] ^ layer_0[669]; 
    assign out[358] = layer_0[131] ^ layer_0[1219]; 
    assign out[359] = ~layer_0[2433]; 
    assign out[360] = layer_0[2352] ^ layer_0[1722]; 
    assign out[361] = ~(layer_0[989] & layer_0[234]); 
    assign out[362] = layer_0[1886] ^ layer_0[574]; 
    assign out[363] = ~layer_0[312] | (layer_0[698] & layer_0[312]); 
    assign out[364] = ~(layer_0[632] & layer_0[2100]); 
    assign out[365] = ~(layer_0[944] & layer_0[421]); 
    assign out[366] = layer_0[132] | layer_0[163]; 
    assign out[367] = ~layer_0[2393] | (layer_0[2301] & layer_0[2393]); 
    assign out[368] = layer_0[1850] ^ layer_0[2297]; 
    assign out[369] = layer_0[2431] ^ layer_0[2309]; 
    assign out[370] = ~(layer_0[1812] ^ layer_0[2513]); 
    assign out[371] = ~(layer_0[1315] ^ layer_0[324]); 
    assign out[372] = ~(layer_0[2108] ^ layer_0[1989]); 
    assign out[373] = layer_0[481]; 
    assign out[374] = ~layer_0[380] | (layer_0[380] & layer_0[938]); 
    assign out[375] = ~(layer_0[704] ^ layer_0[2417]); 
    assign out[376] = ~(layer_0[53] ^ layer_0[412]); 
    assign out[377] = layer_0[617] ^ layer_0[1143]; 
    assign out[378] = ~(layer_0[1895] ^ layer_0[2447]); 
    assign out[379] = layer_0[2325] ^ layer_0[779]; 
    assign out[380] = layer_0[2394] ^ layer_0[2083]; 
    assign out[381] = layer_0[866] ^ layer_0[2049]; 
    assign out[382] = layer_0[362]; 
    assign out[383] = layer_0[1785]; 
    assign out[384] = layer_0[1043]; 
    assign out[385] = ~layer_0[1047] | (layer_0[482] & layer_0[1047]); 
    assign out[386] = ~(layer_0[476] & layer_0[1601]); 
    assign out[387] = layer_0[339] | layer_0[2354]; 
    assign out[388] = layer_0[1712] & ~layer_0[2024]; 
    assign out[389] = ~layer_0[2211] | (layer_0[1469] & layer_0[2211]); 
    assign out[390] = ~(layer_0[1864] ^ layer_0[33]); 
    assign out[391] = ~(layer_0[479] ^ layer_0[1706]); 
    assign out[392] = ~layer_0[447] | (layer_0[447] & layer_0[154]); 
    assign out[393] = layer_0[314] ^ layer_0[354]; 
    assign out[394] = layer_0[1901]; 
    assign out[395] = ~(layer_0[1285] ^ layer_0[2106]); 
    assign out[396] = ~layer_0[1185]; 
    assign out[397] = ~(layer_0[1191] ^ layer_0[2256]); 
    assign out[398] = layer_0[1872] ^ layer_0[296]; 
    assign out[399] = ~(layer_0[1098] ^ layer_0[334]); 
    assign out[400] = ~(layer_0[2517] ^ layer_0[674]); 
    assign out[401] = ~(layer_0[1615] ^ layer_0[1920]); 
    assign out[402] = layer_0[1820]; 
    assign out[403] = layer_0[1669] ^ layer_0[1413]; 
    assign out[404] = layer_0[565] ^ layer_0[1595]; 
    assign out[405] = layer_0[2212] ^ layer_0[375]; 
    assign out[406] = layer_0[1947] & layer_0[1003]; 
    assign out[407] = ~(layer_0[1680] | layer_0[1016]); 
    assign out[408] = layer_0[802] & ~layer_0[179]; 
    assign out[409] = layer_0[1160]; 
    assign out[410] = ~(layer_0[1833] ^ layer_0[648]); 
    assign out[411] = ~(layer_0[673] ^ layer_0[2536]); 
    assign out[412] = layer_0[2508] & layer_0[904]; 
    assign out[413] = layer_0[1318] & layer_0[1766]; 
    assign out[414] = ~(layer_0[780] ^ layer_0[1035]); 
    assign out[415] = ~layer_0[249]; 
    assign out[416] = layer_0[2082] ^ layer_0[1744]; 
    assign out[417] = layer_0[1467] & layer_0[1568]; 
    assign out[418] = ~(layer_0[1133] | layer_0[2476]); 
    assign out[419] = ~layer_0[773]; 
    assign out[420] = layer_0[2124]; 
    assign out[421] = ~(layer_0[469] & layer_0[1023]); 
    assign out[422] = layer_0[1429] ^ layer_0[414]; 
    assign out[423] = layer_0[521] ^ layer_0[665]; 
    assign out[424] = layer_0[1732] ^ layer_0[735]; 
    assign out[425] = ~layer_0[753] | (layer_0[753] & layer_0[1553]); 
    assign out[426] = layer_0[439]; 
    assign out[427] = ~layer_0[1887]; 
    assign out[428] = ~layer_0[1611]; 
    assign out[429] = layer_0[150] & ~layer_0[595]; 
    assign out[430] = layer_0[2080] | layer_0[699]; 
    assign out[431] = ~(layer_0[2298] | layer_0[480]); 
    assign out[432] = ~(layer_0[2037] ^ layer_0[212]); 
    assign out[433] = ~(layer_0[2457] ^ layer_0[534]); 
    assign out[434] = layer_0[2150]; 
    assign out[435] = layer_0[1725]; 
    assign out[436] = layer_0[835] & ~layer_0[405]; 
    assign out[437] = ~layer_0[1907] | (layer_0[1907] & layer_0[1283]); 
    assign out[438] = layer_0[661] ^ layer_0[1423]; 
    assign out[439] = layer_0[2003] ^ layer_0[1985]; 
    assign out[440] = layer_0[2113] & layer_0[994]; 
    assign out[441] = layer_0[2071] | layer_0[1893]; 
    assign out[442] = layer_0[115] ^ layer_0[1343]; 
    assign out[443] = ~layer_0[1193] | (layer_0[610] & layer_0[1193]); 
    assign out[444] = ~(layer_0[1000] & layer_0[2267]); 
    assign out[445] = layer_0[94] ^ layer_0[2273]; 
    assign out[446] = ~(layer_0[1266] ^ layer_0[0]); 
    assign out[447] = layer_0[1777]; 
    assign out[448] = ~layer_0[1264]; 
    assign out[449] = layer_0[505]; 
    assign out[450] = layer_0[877] ^ layer_0[1578]; 
    assign out[451] = ~layer_0[654] | (layer_0[239] & layer_0[654]); 
    assign out[452] = layer_0[2146] & ~layer_0[2209]; 
    assign out[453] = layer_0[201]; 
    assign out[454] = ~(layer_0[162] ^ layer_0[963]); 
    assign out[455] = layer_0[1773]; 
    assign out[456] = layer_0[1376] & ~layer_0[2182]; 
    assign out[457] = ~(layer_0[2554] | layer_0[760]); 
    assign out[458] = ~(layer_0[951] ^ layer_0[408]); 
    assign out[459] = ~layer_0[865] | (layer_0[865] & layer_0[1819]); 
    assign out[460] = layer_0[57] ^ layer_0[2225]; 
    assign out[461] = layer_0[1801] ^ layer_0[633]; 
    assign out[462] = layer_0[2018]; 
    assign out[463] = ~(layer_0[803] ^ layer_0[1771]); 
    assign out[464] = layer_0[1623] & layer_0[2027]; 
    assign out[465] = layer_0[1260] ^ layer_0[1259]; 
    assign out[466] = layer_0[1269]; 
    assign out[467] = ~(layer_0[958] | layer_0[2420]); 
    assign out[468] = layer_0[2528] & ~layer_0[532]; 
    assign out[469] = ~(layer_0[11] ^ layer_0[2034]); 
    assign out[470] = ~(layer_0[465] ^ layer_0[7]); 
    assign out[471] = ~(layer_0[1172] ^ layer_0[1419]); 
    assign out[472] = ~(layer_0[713] ^ layer_0[430]); 
    assign out[473] = ~layer_0[625]; 
    assign out[474] = layer_0[2248]; 
    assign out[475] = layer_0[2230]; 
    assign out[476] = layer_0[454]; 
    assign out[477] = ~(layer_0[1729] | layer_0[942]); 
    assign out[478] = layer_0[689]; 
    assign out[479] = layer_0[543] ^ layer_0[119]; 
    assign out[480] = layer_0[611]; 
    assign out[481] = ~(layer_0[701] ^ layer_0[403]); 
    assign out[482] = ~layer_0[719]; 
    assign out[483] = layer_0[31]; 
    assign out[484] = layer_0[73] & ~layer_0[310]; 
    assign out[485] = ~(layer_0[2556] ^ layer_0[1938]); 
    assign out[486] = ~(layer_0[995] ^ layer_0[1076]); 
    assign out[487] = layer_0[1768] ^ layer_0[2327]; 
    assign out[488] = layer_0[668] ^ layer_0[1758]; 
    assign out[489] = ~(layer_0[614] & layer_0[710]); 
    assign out[490] = ~(layer_0[1439] ^ layer_0[1823]); 
    assign out[491] = ~(layer_0[39] | layer_0[2330]); 
    assign out[492] = ~layer_0[443] | (layer_0[1876] & layer_0[443]); 
    assign out[493] = ~layer_0[427]; 
    assign out[494] = ~layer_0[1711] | (layer_0[1711] & layer_0[1013]); 
    assign out[495] = layer_0[2414] & layer_0[560]; 
    assign out[496] = layer_0[2520] ^ layer_0[464]; 
    assign out[497] = layer_0[1346] & ~layer_0[754]; 
    assign out[498] = ~(layer_0[914] | layer_0[224]); 
    assign out[499] = layer_0[2499]; 
    assign out[500] = layer_0[1742]; 
    assign out[501] = ~layer_0[873] | (layer_0[873] & layer_0[2200]); 
    assign out[502] = layer_0[133]; 
    assign out[503] = ~layer_0[1923] | (layer_0[1923] & layer_0[2466]); 
    assign out[504] = ~(layer_0[554] ^ layer_0[1664]); 
    assign out[505] = layer_0[1821] | layer_0[2126]; 
    assign out[506] = ~layer_0[782]; 
    assign out[507] = ~(layer_0[1239] ^ layer_0[190]); 
    assign out[508] = ~(layer_0[348] ^ layer_0[453]); 
    assign out[509] = layer_0[566] ^ layer_0[723]; 
    assign out[510] = ~(layer_0[1099] & layer_0[1478]); 
    assign out[511] = ~(layer_0[1192] ^ layer_0[736]); 
    assign out[512] = layer_0[1388] & ~layer_0[1404]; 
    assign out[513] = ~layer_0[381]; 
    assign out[514] = layer_0[1500] & layer_0[2347]; 
    assign out[515] = ~layer_0[1916]; 
    assign out[516] = layer_0[1784] & layer_0[600]; 
    assign out[517] = layer_0[2496] & ~layer_0[236]; 
    assign out[518] = layer_0[419] ^ layer_0[607]; 
    assign out[519] = ~(layer_0[207] ^ layer_0[892]); 
    assign out[520] = layer_0[1699] ^ layer_0[1684]; 
    assign out[521] = ~layer_0[594]; 
    assign out[522] = layer_0[2059]; 
    assign out[523] = layer_0[2322]; 
    assign out[524] = layer_0[1097] ^ layer_0[393]; 
    assign out[525] = ~(layer_0[626] ^ layer_0[1406]); 
    assign out[526] = layer_0[886] | layer_0[1021]; 
    assign out[527] = ~layer_0[462]; 
    assign out[528] = ~(layer_0[905] ^ layer_0[693]); 
    assign out[529] = ~(layer_0[1119] | layer_0[1444]); 
    assign out[530] = layer_0[913] ^ layer_0[213]; 
    assign out[531] = ~layer_0[1241] | (layer_0[364] & layer_0[1241]); 
    assign out[532] = ~layer_0[319] | (layer_0[2096] & layer_0[319]); 
    assign out[533] = layer_0[2249]; 
    assign out[534] = layer_0[1797] ^ layer_0[520]; 
    assign out[535] = ~layer_0[1813] | (layer_0[2539] & layer_0[1813]); 
    assign out[536] = ~(layer_0[917] ^ layer_0[1238]); 
    assign out[537] = layer_0[407]; 
    assign out[538] = layer_0[2252] & layer_0[436]; 
    assign out[539] = layer_0[2346]; 
    assign out[540] = layer_0[703] | layer_0[2075]; 
    assign out[541] = ~layer_0[2548]; 
    assign out[542] = layer_0[304] ^ layer_0[2341]; 
    assign out[543] = layer_0[352] ^ layer_0[2235]; 
    assign out[544] = layer_0[2386] ^ layer_0[235]; 
    assign out[545] = layer_0[2540] & ~layer_0[2188]; 
    assign out[546] = layer_0[2253] ^ layer_0[1878]; 
    assign out[547] = ~layer_0[1617]; 
    assign out[548] = ~layer_0[1457]; 
    assign out[549] = ~layer_0[2178] | (layer_0[606] & layer_0[2178]); 
    assign out[550] = layer_0[2236]; 
    assign out[551] = ~layer_0[1027] | (layer_0[1027] & layer_0[923]); 
    assign out[552] = layer_0[1132] ^ layer_0[30]; 
    assign out[553] = ~(layer_0[768] ^ layer_0[1324]); 
    assign out[554] = layer_0[2320] & ~layer_0[316]; 
    assign out[555] = ~layer_0[1182]; 
    assign out[556] = layer_0[1330] & ~layer_0[818]; 
    assign out[557] = ~layer_0[1904]; 
    assign out[558] = layer_0[1188]; 
    assign out[559] = layer_0[1856] ^ layer_0[2455]; 
    assign out[560] = ~(layer_0[1674] ^ layer_0[2224]); 
    assign out[561] = layer_0[1418] ^ layer_0[1361]; 
    assign out[562] = layer_0[511]; 
    assign out[563] = layer_0[712]; 
    assign out[564] = layer_0[240]; 
    assign out[565] = ~layer_0[2276] | (layer_0[2045] & layer_0[2276]); 
    assign out[566] = ~layer_0[1965]; 
    assign out[567] = layer_0[2137] & ~layer_0[1898]; 
    assign out[568] = ~(layer_0[2177] & layer_0[130]); 
    assign out[569] = layer_0[1981] ^ layer_0[2161]; 
    assign out[570] = layer_0[2129]; 
    assign out[571] = layer_0[1978] ^ layer_0[1884]; 
    assign out[572] = layer_0[933] & layer_0[2092]; 
    assign out[573] = layer_0[920] & ~layer_0[714]; 
    assign out[574] = layer_0[1762] ^ layer_0[1905]; 
    assign out[575] = layer_0[874]; 
    assign out[576] = layer_0[2192] & layer_0[70]; 
    assign out[577] = ~layer_0[599]; 
    assign out[578] = layer_0[359]; 
    assign out[579] = layer_0[1533] & layer_0[2522]; 
    assign out[580] = layer_0[2207] & ~layer_0[1869]; 
    assign out[581] = layer_0[1932] ^ layer_0[2110]; 
    assign out[582] = layer_0[158] ^ layer_0[2156]; 
    assign out[583] = layer_0[584]; 
    assign out[584] = layer_0[280] & ~layer_0[848]; 
    assign out[585] = layer_0[623]; 
    assign out[586] = ~(layer_0[27] ^ layer_0[1101]); 
    assign out[587] = layer_0[1689] ^ layer_0[1355]; 
    assign out[588] = layer_0[1695] & ~layer_0[2388]; 
    assign out[589] = layer_0[1633]; 
    assign out[590] = layer_0[1843]; 
    assign out[591] = ~layer_0[2008]; 
    assign out[592] = layer_0[433]; 
    assign out[593] = layer_0[2090] ^ layer_0[1562]; 
    assign out[594] = layer_0[2222] ^ layer_0[613]; 
    assign out[595] = layer_0[2305] | layer_0[897]; 
    assign out[596] = ~(layer_0[1240] ^ layer_0[1325]); 
    assign out[597] = layer_0[747] & ~layer_0[1659]; 
    assign out[598] = layer_0[177] ^ layer_0[1305]; 
    assign out[599] = ~layer_0[425]; 
    assign out[600] = layer_0[898]; 
    assign out[601] = layer_0[587] ^ layer_0[820]; 
    assign out[602] = layer_0[1136] ^ layer_0[2173]; 
    assign out[603] = ~(layer_0[1569] ^ layer_0[1049]); 
    assign out[604] = ~layer_0[2407]; 
    assign out[605] = layer_0[853] & layer_0[470]; 
    assign out[606] = ~(layer_0[1838] | layer_0[2451]); 
    assign out[607] = layer_0[739]; 
    assign out[608] = ~(layer_0[2217] ^ layer_0[2364]); 
    assign out[609] = layer_0[1892]; 
    assign out[610] = layer_0[1628]; 
    assign out[611] = ~(layer_0[1632] ^ layer_0[2530]); 
    assign out[612] = ~layer_0[2390]; 
    assign out[613] = ~layer_0[1782]; 
    assign out[614] = ~layer_0[298]; 
    assign out[615] = layer_0[1105] & ~layer_0[1165]; 
    assign out[616] = layer_0[941]; 
    assign out[617] = layer_0[333] & ~layer_0[690]; 
    assign out[618] = layer_0[1054] | layer_0[896]; 
    assign out[619] = layer_0[2485]; 
    assign out[620] = ~layer_0[2237]; 
    assign out[621] = layer_0[208] & layer_0[242]; 
    assign out[622] = layer_0[385] & ~layer_0[1]; 
    assign out[623] = layer_0[206] ^ layer_0[120]; 
    assign out[624] = layer_0[1311] ^ layer_0[2030]; 
    assign out[625] = layer_0[1026] & ~layer_0[1666]; 
    assign out[626] = layer_0[1248] ^ layer_0[522]; 
    assign out[627] = ~layer_0[544] | (layer_0[544] & layer_0[925]); 
    assign out[628] = ~layer_0[2223] | (layer_0[284] & layer_0[2223]); 
    assign out[629] = ~(layer_0[74] ^ layer_0[2509]); 
    assign out[630] = layer_0[347] & layer_0[2012]; 
    assign out[631] = layer_0[248] ^ layer_0[1494]; 
    assign out[632] = layer_0[2153] ^ layer_0[2488]; 
    assign out[633] = layer_0[1804] & layer_0[1922]; 
    assign out[634] = layer_0[1431]; 
    assign out[635] = ~layer_0[92]; 
    assign out[636] = layer_0[979]; 
    assign out[637] = layer_0[720] ^ layer_0[1882]; 
    assign out[638] = ~(layer_0[801] | layer_0[1358]); 
    assign out[639] = layer_0[1506] & ~layer_0[2149]; 
    assign out[640] = ~(layer_0[858] ^ layer_0[129]); 
    assign out[641] = ~(layer_0[1509] ^ layer_0[1523]); 
    assign out[642] = ~(layer_0[200] & layer_0[1225]); 
    assign out[643] = layer_0[851] ^ layer_0[1501]; 
    assign out[644] = layer_0[1381]; 
    assign out[645] = layer_0[1842] ^ layer_0[1673]; 
    assign out[646] = ~layer_0[281] | (layer_0[1903] & layer_0[281]); 
    assign out[647] = ~(layer_0[99] ^ layer_0[1137]); 
    assign out[648] = layer_0[1492]; 
    assign out[649] = ~(layer_0[1860] ^ layer_0[965]); 
    assign out[650] = ~layer_0[1111]; 
    assign out[651] = layer_0[2020]; 
    assign out[652] = ~layer_0[2218]; 
    assign out[653] = layer_0[2316] ^ layer_0[285]; 
    assign out[654] = ~layer_0[1504]; 
    assign out[655] = ~layer_0[1073] | (layer_0[1399] & layer_0[1073]); 
    assign out[656] = ~(layer_0[1924] ^ layer_0[2041]); 
    assign out[657] = layer_0[927] ^ layer_0[1848]; 
    assign out[658] = ~layer_0[2337]; 
    assign out[659] = layer_0[2400] ^ layer_0[2521]; 
    assign out[660] = ~layer_0[58]; 
    assign out[661] = layer_0[1958] ^ layer_0[809]; 
    assign out[662] = ~(layer_0[320] ^ layer_0[2446]); 
    assign out[663] = ~(layer_0[1670] | layer_0[928]); 
    assign out[664] = ~(layer_0[1433] ^ layer_0[1557]); 
    assign out[665] = layer_0[328] | layer_0[1279]; 
    assign out[666] = layer_0[1256] & ~layer_0[1675]; 
    assign out[667] = layer_0[1234] ^ layer_0[663]; 
    assign out[668] = layer_0[2434] ^ layer_0[664]; 
    assign out[669] = layer_0[1396] & ~layer_0[1906]; 
    assign out[670] = layer_0[2238] | layer_0[696]; 
    assign out[671] = layer_0[1454] ^ layer_0[1941]; 
    assign out[672] = ~(layer_0[437] | layer_0[1542]); 
    assign out[673] = ~layer_0[1832]; 
    assign out[674] = layer_0[1100] | layer_0[1180]; 
    assign out[675] = ~(layer_0[434] ^ layer_0[1432]); 
    assign out[676] = layer_0[855] ^ layer_0[2133]; 
    assign out[677] = layer_0[1373] ^ layer_0[1150]; 
    assign out[678] = ~(layer_0[1873] ^ layer_0[812]); 
    assign out[679] = layer_0[1018] ^ layer_0[1201]; 
    assign out[680] = ~layer_0[1448] | (layer_0[1448] & layer_0[1139]); 
    assign out[681] = layer_0[564] ^ layer_0[124]; 
    assign out[682] = layer_0[980]; 
    assign out[683] = layer_0[2140] ^ layer_0[466]; 
    assign out[684] = layer_0[2399] & ~layer_0[1942]; 
    assign out[685] = ~layer_0[1716] | (layer_0[1752] & layer_0[1716]); 
    assign out[686] = ~(layer_0[1218] & layer_0[1663]); 
    assign out[687] = layer_0[88] ^ layer_0[1287]; 
    assign out[688] = layer_0[2219]; 
    assign out[689] = ~layer_0[8] | (layer_0[8] & layer_0[738]); 
    assign out[690] = ~layer_0[749]; 
    assign out[691] = layer_0[93] | layer_0[452]; 
    assign out[692] = ~(layer_0[61] & layer_0[1345]); 
    assign out[693] = ~layer_0[725] | (layer_0[2125] & layer_0[725]); 
    assign out[694] = ~layer_0[199] | (layer_0[199] & layer_0[1583]); 
    assign out[695] = ~layer_0[1295]; 
    assign out[696] = ~(layer_0[881] ^ layer_0[581]); 
    assign out[697] = layer_0[1371]; 
    assign out[698] = layer_0[2366] | layer_0[901]; 
    assign out[699] = layer_0[241]; 
    assign out[700] = layer_0[1383] & ~layer_0[180]; 
    assign out[701] = ~(layer_0[539] ^ layer_0[170]); 
    assign out[702] = layer_0[1528] & layer_0[2290]; 
    assign out[703] = layer_0[1621]; 
    assign out[704] = layer_0[2170] ^ layer_0[680]; 
    assign out[705] = layer_0[1207] & ~layer_0[151]; 
    assign out[706] = layer_0[1622]; 
    assign out[707] = layer_0[459] ^ layer_0[378]; 
    assign out[708] = layer_0[1900] | layer_0[72]; 
    assign out[709] = layer_0[2487] | layer_0[397]; 
    assign out[710] = layer_0[467] ^ layer_0[220]; 
    assign out[711] = ~layer_0[127]; 
    assign out[712] = layer_0[1299] ^ layer_0[1915]; 
    assign out[713] = layer_0[570] ^ layer_0[509]; 
    assign out[714] = layer_0[640] ^ layer_0[114]; 
    assign out[715] = ~layer_0[1713]; 
    assign out[716] = ~(layer_0[1626] ^ layer_0[3]); 
    assign out[717] = layer_0[2537]; 
    assign out[718] = layer_0[2461]; 
    assign out[719] = layer_0[656] & ~layer_0[597]; 
    assign out[720] = layer_0[1007] | layer_0[2445]; 
    assign out[721] = layer_0[1890] & ~layer_0[2524]; 
    assign out[722] = layer_0[862]; 
    assign out[723] = ~layer_0[2231]; 
    assign out[724] = ~(layer_0[1983] | layer_0[1110]); 
    assign out[725] = ~(layer_0[76] ^ layer_0[2077]); 
    assign out[726] = layer_0[2138]; 
    assign out[727] = layer_0[100]; 
    assign out[728] = layer_0[157]; 
    assign out[729] = layer_0[1827] | layer_0[1233]; 
    assign out[730] = ~(layer_0[1216] ^ layer_0[184]); 
    assign out[731] = layer_0[13] | layer_0[1147]; 
    assign out[732] = ~layer_0[2042] | (layer_0[1118] & layer_0[2042]); 
    assign out[733] = layer_0[2085]; 
    assign out[734] = layer_0[1322]; 
    assign out[735] = layer_0[20]; 
    assign out[736] = layer_0[1462]; 
    assign out[737] = ~layer_0[628]; 
    assign out[738] = layer_0[2419] | layer_0[118]; 
    assign out[739] = layer_0[798] ^ layer_0[139]; 
    assign out[740] = layer_0[2356] | layer_0[970]; 
    assign out[741] = ~layer_0[2065]; 
    assign out[742] = layer_0[410] ^ layer_0[879]; 
    assign out[743] = layer_0[2016] ^ layer_0[1296]; 
    assign out[744] = layer_0[2275] ^ layer_0[1954]; 
    assign out[745] = ~(layer_0[919] ^ layer_0[612]); 
    assign out[746] = ~layer_0[1921]; 
    assign out[747] = layer_0[1142] | layer_0[1113]; 
    assign out[748] = layer_0[1340] & layer_0[1585]; 
    assign out[749] = layer_0[18] & layer_0[1434]; 
    assign out[750] = layer_0[2492]; 
    assign out[751] = ~layer_0[1547]; 
    assign out[752] = layer_0[1080] & layer_0[847]; 
    assign out[753] = layer_0[321]; 
    assign out[754] = layer_0[1556] ^ layer_0[1751]; 
    assign out[755] = layer_0[1129] ^ layer_0[1391]; 
    assign out[756] = layer_0[526] & layer_0[2169]; 
    assign out[757] = layer_0[2323] & ~layer_0[1963]; 
    assign out[758] = ~(layer_0[2265] ^ layer_0[1554]); 
    assign out[759] = layer_0[1704] | layer_0[2378]; 
    assign out[760] = ~(layer_0[1057] ^ layer_0[1470]); 
    assign out[761] = layer_0[1290] | layer_0[440]; 
    assign out[762] = layer_0[1055] & ~layer_0[1787]; 
    assign out[763] = ~layer_0[1959]; 
    assign out[764] = layer_0[745] ^ layer_0[261]; 
    assign out[765] = ~(layer_0[493] & layer_0[2262]); 
    assign out[766] = layer_0[2141] & ~layer_0[1849]; 
    assign out[767] = layer_0[2438] ^ layer_0[1815]; 
    assign out[768] = ~(layer_0[1576] ^ layer_0[953]); 
    assign out[769] = ~layer_0[691]; 
    assign out[770] = layer_0[2198] ^ layer_0[2481]; 
    assign out[771] = ~layer_0[1117]; 
    assign out[772] = layer_0[2334] ^ layer_0[1032]; 
    assign out[773] = layer_0[2437] ^ layer_0[685]; 
    assign out[774] = ~(layer_0[2348] | layer_0[1366]); 
    assign out[775] = layer_0[1034]; 
    assign out[776] = layer_0[1580] ^ layer_0[637]; 
    assign out[777] = layer_0[1960] ^ layer_0[1846]; 
    assign out[778] = layer_0[1029] & ~layer_0[1988]; 
    assign out[779] = layer_0[921] & ~layer_0[1612]; 
    assign out[780] = layer_0[1607] & ~layer_0[646]; 
    assign out[781] = ~(layer_0[1417] & layer_0[416]); 
    assign out[782] = ~(layer_0[1514] & layer_0[1507]); 
    assign out[783] = ~(layer_0[967] | layer_0[2436]); 
    assign out[784] = ~(layer_0[1714] | layer_0[2116]); 
    assign out[785] = layer_0[1354] & ~layer_0[1255]; 
    assign out[786] = layer_0[1041] & ~layer_0[1227]; 
    assign out[787] = layer_0[863] | layer_0[149]; 
    assign out[788] = ~layer_0[732]; 
    assign out[789] = layer_0[2164] & ~layer_0[370]; 
    assign out[790] = layer_0[791] & ~layer_0[1177]; 
    assign out[791] = layer_0[2515] & layer_0[2470]; 
    assign out[792] = ~layer_0[533] | (layer_0[533] & layer_0[116]); 
    assign out[793] = layer_0[1571] & ~layer_0[489]; 
    assign out[794] = layer_0[592] & ~layer_0[1912]; 
    assign out[795] = ~layer_0[1485] | (layer_0[1385] & layer_0[1485]); 
    assign out[796] = layer_0[2359] & layer_0[203]; 
    assign out[797] = layer_0[887]; 
    assign out[798] = ~layer_0[514]; 
    assign out[799] = ~(layer_0[1070] ^ layer_0[961]); 
    assign out[800] = layer_0[2353] & ~layer_0[1116]; 
    assign out[801] = ~(layer_0[804] | layer_0[1756]); 
    assign out[802] = layer_0[645] ^ layer_0[1449]; 
    assign out[803] = layer_0[490] ^ layer_0[2208]; 
    assign out[804] = ~layer_0[2168]; 
    assign out[805] = layer_0[501] & ~layer_0[1949]; 
    assign out[806] = ~(layer_0[785] ^ layer_0[2312]); 
    assign out[807] = layer_0[678] & layer_0[1519]; 
    assign out[808] = ~layer_0[2396]; 
    assign out[809] = ~(layer_0[2098] | layer_0[1088]); 
    assign out[810] = layer_0[1979] & layer_0[755]; 
    assign out[811] = layer_0[2529] ^ layer_0[2254]; 
    assign out[812] = layer_0[1228] ^ layer_0[2115]; 
    assign out[813] = ~(layer_0[2000] ^ layer_0[1422]); 
    assign out[814] = ~(layer_0[1908] | layer_0[2454]); 
    assign out[815] = ~layer_0[161]; 
    assign out[816] = layer_0[997] & ~layer_0[1505]; 
    assign out[817] = ~layer_0[1208]; 
    assign out[818] = layer_0[125] & layer_0[1199]; 
    assign out[819] = layer_0[1593] & ~layer_0[1527]; 
    assign out[820] = layer_0[89] & ~layer_0[1997]; 
    assign out[821] = layer_0[483] & ~layer_0[830]; 
    assign out[822] = layer_0[2191] & layer_0[695]; 
    assign out[823] = ~(layer_0[1254] ^ layer_0[1943]); 
    assign out[824] = ~layer_0[2004] | (layer_0[528] & layer_0[2004]); 
    assign out[825] = ~layer_0[1871] | (layer_0[1871] & layer_0[289]); 
    assign out[826] = layer_0[288] ^ layer_0[702]; 
    assign out[827] = layer_0[596] ^ layer_0[1745]; 
    assign out[828] = layer_0[143]; 
    assign out[829] = layer_0[2180] & ~layer_0[1982]; 
    assign out[830] = ~layer_0[1753]; 
    assign out[831] = layer_0[583] & layer_0[1564]; 
    assign out[832] = ~(layer_0[1735] ^ layer_0[1570]); 
    assign out[833] = layer_0[900]; 
    assign out[834] = layer_0[2111] ^ layer_0[223]; 
    assign out[835] = ~(layer_0[513] | layer_0[605]); 
    assign out[836] = ~(layer_0[1427] | layer_0[1881]); 
    assign out[837] = layer_0[1006] | layer_0[1661]; 
    assign out[838] = ~(layer_0[2291] ^ layer_0[176]); 
    assign out[839] = ~(layer_0[1465] ^ layer_0[1438]); 
    assign out[840] = ~layer_0[451]; 
    assign out[841] = ~(layer_0[2443] | layer_0[2233]); 
    assign out[842] = layer_0[1624] & layer_0[1754]; 
    assign out[843] = layer_0[2439] ^ layer_0[2373]; 
    assign out[844] = layer_0[1831] & ~layer_0[2009]; 
    assign out[845] = ~(layer_0[1640] ^ layer_0[1186]); 
    assign out[846] = layer_0[1822] & ~layer_0[2377]; 
    assign out[847] = layer_0[2313] & ~layer_0[655]; 
    assign out[848] = layer_0[2] & ~layer_0[1171]; 
    assign out[849] = ~(layer_0[2176] & layer_0[315]); 
    assign out[850] = layer_0[1521] & ~layer_0[2507]; 
    assign out[851] = ~layer_0[946]; 
    assign out[852] = layer_0[1854]; 
    assign out[853] = layer_0[1529] & ~layer_0[1362]; 
    assign out[854] = layer_0[43]; 
    assign out[855] = ~layer_0[1202]; 
    assign out[856] = layer_0[1493] ^ layer_0[2463]; 
    assign out[857] = layer_0[2272] ^ layer_0[1934]; 
    assign out[858] = ~layer_0[428]; 
    assign out[859] = layer_0[204] & ~layer_0[394]; 
    assign out[860] = ~(layer_0[2401] ^ layer_0[1477]); 
    assign out[861] = layer_0[1718] ^ layer_0[1048]; 
    assign out[862] = ~layer_0[1910] | (layer_0[1534] & layer_0[1910]); 
    assign out[863] = layer_0[2478]; 
    assign out[864] = ~(layer_0[2143] ^ layer_0[349]); 
    assign out[865] = layer_0[384] | layer_0[959]; 
    assign out[866] = layer_0[2058] & layer_0[1144]; 
    assign out[867] = ~(layer_0[2278] ^ layer_0[1840]); 
    assign out[868] = ~layer_0[1377] | (layer_0[639] & layer_0[1377]); 
    assign out[869] = ~(layer_0[1309] ^ layer_0[1894]); 
    assign out[870] = ~layer_0[590]; 
    assign out[871] = layer_0[650] & ~layer_0[1342]; 
    assign out[872] = ~layer_0[142] | (layer_0[142] & layer_0[1044]); 
    assign out[873] = ~layer_0[269] | (layer_0[1151] & layer_0[269]); 
    assign out[874] = layer_0[758] & ~layer_0[984]; 
    assign out[875] = layer_0[1733] ^ layer_0[1897]; 
    assign out[876] = ~layer_0[471]; 
    assign out[877] = layer_0[2121] & layer_0[1360]; 
    assign out[878] = ~(layer_0[842] ^ layer_0[1440]); 
    assign out[879] = layer_0[1223] & layer_0[1247]; 
    assign out[880] = layer_0[1014]; 
    assign out[881] = layer_0[1083]; 
    assign out[882] = ~(layer_0[1613] ^ layer_0[2199]); 
    assign out[883] = layer_0[257]; 
    assign out[884] = layer_0[1654] | layer_0[1039]; 
    assign out[885] = layer_0[1579] | layer_0[2306]; 
    assign out[886] = ~(layer_0[376] ^ layer_0[722]); 
    assign out[887] = ~layer_0[1235]; 
    assign out[888] = layer_0[1224] & ~layer_0[2295]; 
    assign out[889] = ~(layer_0[95] ^ layer_0[1721]); 
    assign out[890] = ~layer_0[263]; 
    assign out[891] = layer_0[567] & layer_0[1510]; 
    assign out[892] = ~layer_0[1442] | (layer_0[2398] & layer_0[1442]); 
    assign out[893] = layer_0[2489] & ~layer_0[1271]; 
    assign out[894] = ~layer_0[1880]; 
    assign out[895] = ~layer_0[795]; 
    assign out[896] = layer_0[2010] & ~layer_0[2119]; 
    assign out[897] = layer_0[519] ^ layer_0[1495]; 
    assign out[898] = ~(layer_0[1925] ^ layer_0[1750]); 
    assign out[899] = layer_0[1852] & layer_0[49]; 
    assign out[900] = layer_0[1676] ^ layer_0[1660]; 
    assign out[901] = ~layer_0[759]; 
    assign out[902] = layer_0[1334] ^ layer_0[2193]; 
    assign out[903] = layer_0[1336]; 
    assign out[904] = layer_0[1268] & ~layer_0[1437]; 
    assign out[905] = layer_0[387] & ~layer_0[2532]; 
    assign out[906] = ~layer_0[1230]; 
    assign out[907] = layer_0[2404] ^ layer_0[867]; 
    assign out[908] = ~(layer_0[692] & layer_0[1575]); 
    assign out[909] = ~(layer_0[463] | layer_0[1486]); 
    assign out[910] = ~(layer_0[1480] ^ layer_0[1456]); 
    assign out[911] = ~layer_0[2268] | (layer_0[2268] & layer_0[2360]); 
    assign out[912] = layer_0[307] | layer_0[2118]; 
    assign out[913] = layer_0[2094] & layer_0[1555]; 
    assign out[914] = layer_0[1320] & ~layer_0[1550]; 
    assign out[915] = layer_0[1002] & layer_0[2333]; 
    assign out[916] = layer_0[1788] & ~layer_0[1630]; 
    assign out[917] = ~(layer_0[2501] | layer_0[990]); 
    assign out[918] = layer_0[1899] & layer_0[1265]; 
    assign out[919] = ~(layer_0[1169] ^ layer_0[84]); 
    assign out[920] = layer_0[1642]; 
    assign out[921] = layer_0[744] | layer_0[1019]; 
    assign out[922] = layer_0[2175] & ~layer_0[1036]; 
    assign out[923] = layer_0[604] & ~layer_0[864]; 
    assign out[924] = ~layer_0[2541]; 
    assign out[925] = layer_0[2220] ^ layer_0[1168]; 
    assign out[926] = ~(layer_0[1213] ^ layer_0[2319]); 
    assign out[927] = layer_0[1069] ^ layer_0[2289]; 
    assign out[928] = ~(layer_0[884] | layer_0[2480]); 
    assign out[929] = layer_0[1078] ^ layer_0[844]; 
    assign out[930] = ~(layer_0[662] | layer_0[1599]); 
    assign out[931] = layer_0[1331] & layer_0[1602]; 
    assign out[932] = layer_0[789] & layer_0[2300]; 
    assign out[933] = ~(layer_0[1865] ^ layer_0[1896]); 
    assign out[934] = ~(layer_0[1491] ^ layer_0[305]); 
    assign out[935] = ~layer_0[2073]; 
    assign out[936] = ~(layer_0[2165] | layer_0[2387]); 
    assign out[937] = layer_0[360]; 
    assign out[938] = layer_0[1902] & layer_0[1760]; 
    assign out[939] = ~(layer_0[841] ^ layer_0[1929]); 
    assign out[940] = ~(layer_0[978] | layer_0[2435]); 
    assign out[941] = layer_0[311]; 
    assign out[942] = ~(layer_0[907] | layer_0[2120]); 
    assign out[943] = layer_0[1061]; 
    assign out[944] = ~(layer_0[1148] ^ layer_0[172]); 
    assign out[945] = ~layer_0[2017]; 
    assign out[946] = layer_0[1844] | layer_0[1563]; 
    assign out[947] = layer_0[2117] & ~layer_0[396]; 
    assign out[948] = layer_0[10] & ~layer_0[2338]; 
    assign out[949] = ~(layer_0[1875] | layer_0[247]); 
    assign out[950] = ~(layer_0[618] ^ layer_0[2194]); 
    assign out[951] = ~layer_0[442] | (layer_0[367] & layer_0[442]); 
    assign out[952] = ~(layer_0[2411] ^ layer_0[922]); 
    assign out[953] = ~layer_0[563]; 
    assign out[954] = ~layer_0[1411]; 
    assign out[955] = layer_0[2385] & layer_0[677]; 
    assign out[956] = layer_0[833] & layer_0[2391]; 
    assign out[957] = layer_0[2091] & layer_0[1962]; 
    assign out[958] = ~layer_0[2244]; 
    assign out[959] = ~(layer_0[1696] ^ layer_0[718]); 
    assign out[960] = ~(layer_0[987] & layer_0[438]); 
    assign out[961] = layer_0[2068] & layer_0[1161]; 
    assign out[962] = layer_0[1928] ^ layer_0[971]; 
    assign out[963] = layer_0[91] ^ layer_0[159]; 
    assign out[964] = layer_0[1763] ^ layer_0[1090]; 
    assign out[965] = layer_0[1022] ^ layer_0[1998]; 
    assign out[966] = ~layer_0[108]; 
    assign out[967] = ~(layer_0[2495] ^ layer_0[392]); 
    assign out[968] = layer_0[1648] ^ layer_0[831]; 
    assign out[969] = ~layer_0[2081] | (layer_0[2081] & layer_0[1122]); 
    assign out[970] = ~(layer_0[1868] | layer_0[2533]); 
    assign out[971] = ~layer_0[1094]; 
    assign out[972] = ~layer_0[1405]; 
    assign out[973] = ~layer_0[2549]; 
    assign out[974] = ~layer_0[1297]; 
    assign out[975] = layer_0[2127] & layer_0[1541]; 
    assign out[976] = layer_0[1891]; 
    assign out[977] = layer_0[2441] & ~layer_0[762]; 
    assign out[978] = ~(layer_0[1879] | layer_0[1679]); 
    assign out[979] = layer_0[110] & layer_0[1747]; 
    assign out[980] = ~(layer_0[2370] ^ layer_0[1244]); 
    assign out[981] = layer_0[889]; 
    assign out[982] = layer_0[1025] & ~layer_0[237]; 
    assign out[983] = layer_0[2050] & ~layer_0[1327]; 
    assign out[984] = layer_0[1987] ^ layer_0[775]; 
    assign out[985] = layer_0[788] & ~layer_0[361]; 
    assign out[986] = ~(layer_0[1079] ^ layer_0[1243]); 
    assign out[987] = layer_0[1977] ^ layer_0[1776]; 
    assign out[988] = layer_0[1306]; 
    assign out[989] = layer_0[1835] | layer_0[2282]; 
    assign out[990] = layer_0[504] & ~layer_0[173]; 
    assign out[991] = ~layer_0[166]; 
    assign out[992] = layer_0[1416] & ~layer_0[1582]; 
    assign out[993] = ~(layer_0[2460] & layer_0[377]); 
    assign out[994] = layer_0[297] & layer_0[1428]; 
    assign out[995] = ~(layer_0[1068] ^ layer_0[629]); 
    assign out[996] = ~layer_0[54]; 
    assign out[997] = layer_0[209]; 
    assign out[998] = layer_0[189] & layer_0[2367]; 
    assign out[999] = layer_0[1293]; 
    assign out[1000] = layer_0[153] & ~layer_0[1765]; 
    assign out[1001] = ~(layer_0[2469] | layer_0[2154]); 
    assign out[1002] = layer_0[420] ^ layer_0[1481]; 
    assign out[1003] = layer_0[2471]; 
    assign out[1004] = layer_0[422] & ~layer_0[191]; 
    assign out[1005] = layer_0[65] & ~layer_0[549]; 
    assign out[1006] = ~(layer_0[659] & layer_0[2304]); 
    assign out[1007] = layer_0[457]; 
    assign out[1008] = ~(layer_0[2221] ^ layer_0[2557]); 
    assign out[1009] = layer_0[1513] & ~layer_0[598]; 
    assign out[1010] = ~layer_0[1638]; 
    assign out[1011] = layer_0[1300]; 
    assign out[1012] = layer_0[323] ^ layer_0[572]; 
    assign out[1013] = layer_0[1598] & layer_0[1359]; 
    assign out[1014] = ~(layer_0[2546] | layer_0[1401]); 
    assign out[1015] = layer_0[1665] ^ layer_0[2060]; 
    assign out[1016] = ~(layer_0[1866] ^ layer_0[2216]); 
    assign out[1017] = ~(layer_0[494] ^ layer_0[1479]); 
    assign out[1018] = layer_0[36]; 
    assign out[1019] = ~layer_0[636]; 
    assign out[1020] = layer_0[426] ^ layer_0[64]; 
    assign out[1021] = ~layer_0[796]; 
    assign out[1022] = layer_0[2122] ^ layer_0[608]; 
    assign out[1023] = ~(layer_0[1253] & layer_0[1531]); 
    assign out[1024] = layer_0[1686] ^ layer_0[2247]; 
    assign out[1025] = layer_0[1056] & layer_0[1559]; 
    assign out[1026] = layer_0[2203] ^ layer_0[1278]; 
    assign out[1027] = ~(layer_0[210] ^ layer_0[1166]); 
    assign out[1028] = ~(layer_0[1141] ^ layer_0[2250]); 
    assign out[1029] = ~(layer_0[939] & layer_0[2344]); 
    assign out[1030] = layer_0[1774] ^ layer_0[546]; 
    assign out[1031] = layer_0[1203] & layer_0[550]; 
    assign out[1032] = ~(layer_0[77] & layer_0[97]); 
    assign out[1033] = layer_0[2181] ^ layer_0[603]; 
    assign out[1034] = ~(layer_0[409] ^ layer_0[1367]); 
    assign out[1035] = ~layer_0[1918]; 
    assign out[1036] = layer_0[609] & layer_0[1772]; 
    assign out[1037] = ~(layer_0[1828] & layer_0[667]); 
    assign out[1038] = ~layer_0[294]; 
    assign out[1039] = ~(layer_0[1275] ^ layer_0[1780]); 
    assign out[1040] = layer_0[337] ^ layer_0[2429]; 
    assign out[1041] = layer_0[40] & ~layer_0[44]; 
    assign out[1042] = ~(layer_0[591] ^ layer_0[1803]); 
    assign out[1043] = layer_0[1280] & ~layer_0[2204]; 
    assign out[1044] = ~(layer_0[1384] ^ layer_0[83]); 
    assign out[1045] = ~(layer_0[1739] ^ layer_0[647]); 
    assign out[1046] = layer_0[500]; 
    assign out[1047] = ~(layer_0[828] ^ layer_0[211]); 
    assign out[1048] = ~(layer_0[278] ^ layer_0[2328]); 
    assign out[1049] = ~(layer_0[2335] ^ layer_0[1786]); 
    assign out[1050] = layer_0[956]; 
    assign out[1051] = ~(layer_0[1525] ^ layer_0[2259]); 
    assign out[1052] = layer_0[1489] ^ layer_0[849]; 
    assign out[1053] = layer_0[1913] & ~layer_0[1112]; 
    assign out[1054] = ~(layer_0[576] ^ layer_0[1955]); 
    assign out[1055] = layer_0[1968] ^ layer_0[822]; 
    assign out[1056] = ~layer_0[63]; 
    assign out[1057] = ~(layer_0[2380] ^ layer_0[2190]); 
    assign out[1058] = layer_0[986] ^ layer_0[1995]; 
    assign out[1059] = ~layer_0[2486] | (layer_0[1692] & layer_0[2486]); 
    assign out[1060] = layer_0[2415]; 
    assign out[1061] = layer_0[1730] ^ layer_0[188]; 
    assign out[1062] = layer_0[2035] ^ layer_0[260]; 
    assign out[1063] = layer_0[98]; 
    assign out[1064] = ~layer_0[1008]; 
    assign out[1065] = ~(layer_0[977] ^ layer_0[1524]); 
    assign out[1066] = layer_0[1859] ^ layer_0[2547]; 
    assign out[1067] = layer_0[774] & layer_0[251]; 
    assign out[1068] = layer_0[1237]; 
    assign out[1069] = ~layer_0[1059]; 
    assign out[1070] = layer_0[1536] ^ layer_0[771]; 
    assign out[1071] = layer_0[411]; 
    assign out[1072] = layer_0[1681]; 
    assign out[1073] = ~layer_0[819] | (layer_0[819] & layer_0[2036]); 
    assign out[1074] = layer_0[1522] & ~layer_0[353]; 
    assign out[1075] = layer_0[834] ^ layer_0[1298]; 
    assign out[1076] = ~(layer_0[1688] ^ layer_0[1028]); 
    assign out[1077] = layer_0[4] | layer_0[1727]; 
    assign out[1078] = ~(layer_0[15] ^ layer_0[2087]); 
    assign out[1079] = layer_0[1351] | layer_0[1154]; 
    assign out[1080] = layer_0[2405] | layer_0[579]; 
    assign out[1081] = layer_0[815] ^ layer_0[1326]; 
    assign out[1082] = ~(layer_0[817] ^ layer_0[460]); 
    assign out[1083] = layer_0[1775] ^ layer_0[2029]; 
    assign out[1084] = layer_0[1370] & layer_0[1066]; 
    assign out[1085] = ~(layer_0[1805] ^ layer_0[25]); 
    assign out[1086] = layer_0[2277] & ~layer_0[2286]; 
    assign out[1087] = layer_0[71]; 
    assign out[1088] = ~layer_0[2032]; 
    assign out[1089] = layer_0[552]; 
    assign out[1090] = layer_0[683] ^ layer_0[2142]; 
    assign out[1091] = ~(layer_0[2038] ^ layer_0[1421]); 
    assign out[1092] = layer_0[756] & ~layer_0[2274]; 
    assign out[1093] = layer_0[1468]; 
    assign out[1094] = ~layer_0[2358]; 
    assign out[1095] = layer_0[455] & layer_0[1526]; 
    assign out[1096] = ~layer_0[733]; 
    assign out[1097] = layer_0[1789] & layer_0[541]; 
    assign out[1098] = layer_0[1252] ^ layer_0[1743]; 
    assign out[1099] = layer_0[631] | layer_0[1231]; 
    assign out[1100] = ~layer_0[1374]; 
    assign out[1101] = ~(layer_0[228] | layer_0[2162]); 
    assign out[1102] = ~layer_0[1045]; 
    assign out[1103] = ~(layer_0[2543] ^ layer_0[1209]); 
    assign out[1104] = layer_0[742]; 
    assign out[1105] = layer_0[1565] ^ layer_0[2475]; 
    assign out[1106] = layer_0[1052] & ~layer_0[331]; 
    assign out[1107] = layer_0[1845]; 
    assign out[1108] = layer_0[823]; 
    assign out[1109] = layer_0[2363] | layer_0[974]; 
    assign out[1110] = layer_0[366]; 
    assign out[1111] = layer_0[2473] & ~layer_0[75]; 
    assign out[1112] = layer_0[1038]; 
    assign out[1113] = layer_0[1667] ^ layer_0[1173]; 
    assign out[1114] = ~(layer_0[168] ^ layer_0[2418]); 
    assign out[1115] = layer_0[906] ^ layer_0[916]; 
    assign out[1116] = ~layer_0[871] | (layer_0[233] & layer_0[871]); 
    assign out[1117] = ~layer_0[1167]; 
    assign out[1118] = layer_0[1198] ^ layer_0[1020]; 
    assign out[1119] = layer_0[113] ^ layer_0[290]; 
    assign out[1120] = ~(layer_0[214] ^ layer_0[498]); 
    assign out[1121] = layer_0[1597] & ~layer_0[2251]; 
    assign out[1122] = ~(layer_0[1826] ^ layer_0[1969]); 
    assign out[1123] = ~layer_0[2206]; 
    assign out[1124] = layer_0[2383] ^ layer_0[535]; 
    assign out[1125] = ~layer_0[503]; 
    assign out[1126] = layer_0[697]; 
    assign out[1127] = ~layer_0[1652] | (layer_0[1652] & layer_0[1811]); 
    assign out[1128] = ~(layer_0[254] ^ layer_0[1096]); 
    assign out[1129] = layer_0[2148] | layer_0[527]; 
    assign out[1130] = ~layer_0[106]; 
    assign out[1131] = layer_0[1120]; 
    assign out[1132] = layer_0[499] & ~layer_0[2023]; 
    assign out[1133] = layer_0[1964]; 
    assign out[1134] = layer_0[1222] ^ layer_0[2351]; 
    assign out[1135] = layer_0[1046] ^ layer_0[2484]; 
    assign out[1136] = layer_0[21] ^ layer_0[1163]; 
    assign out[1137] = ~(layer_0[141] ^ layer_0[1836]); 
    assign out[1138] = ~layer_0[78]; 
    assign out[1139] = ~(layer_0[1138] ^ layer_0[231]); 
    assign out[1140] = ~(layer_0[1135] ^ layer_0[2246]); 
    assign out[1141] = ~(layer_0[1157] ^ layer_0[2232]); 
    assign out[1142] = layer_0[2019] & layer_0[507]; 
    assign out[1143] = layer_0[1459] & ~layer_0[2101]; 
    assign out[1144] = ~(layer_0[1520] ^ layer_0[1512]); 
    assign out[1145] = layer_0[69]; 
    assign out[1146] = layer_0[229] ^ layer_0[777]; 
    assign out[1147] = ~(layer_0[1545] ^ layer_0[2409]); 
    assign out[1148] = layer_0[729] & layer_0[1647]; 
    assign out[1149] = layer_0[1996] ^ layer_0[1037]; 
    assign out[1150] = layer_0[837] & ~layer_0[448]; 
    assign out[1151] = ~(layer_0[1175] | layer_0[1976]); 
    assign out[1152] = ~(layer_0[553] | layer_0[2329]); 
    assign out[1153] = ~(layer_0[1572] ^ layer_0[186]); 
    assign out[1154] = layer_0[80] & layer_0[52]; 
    assign out[1155] = ~(layer_0[1319] | layer_0[2491]); 
    assign out[1156] = layer_0[1511] ^ layer_0[1140]; 
    assign out[1157] = ~(layer_0[2171] | layer_0[562]); 
    assign out[1158] = layer_0[140]; 
    assign out[1159] = layer_0[23] & ~layer_0[1847]; 
    assign out[1160] = layer_0[1728] & ~layer_0[308]; 
    assign out[1161] = layer_0[46] ^ layer_0[1719]; 
    assign out[1162] = ~(layer_0[90] | layer_0[2039]); 
    assign out[1163] = layer_0[2375] & ~layer_0[1292]; 
    assign out[1164] = layer_0[1967]; 
    assign out[1165] = ~(layer_0[955] ^ layer_0[557]); 
    assign out[1166] = ~(layer_0[772] ^ layer_0[356]); 
    assign out[1167] = layer_0[1950] ^ layer_0[2239]; 
    assign out[1168] = ~layer_0[1206]; 
    assign out[1169] = ~(layer_0[136] ^ layer_0[369]); 
    assign out[1170] = layer_0[146] ^ layer_0[2511]; 
    assign out[1171] = ~(layer_0[1220] ^ layer_0[1072]); 
    assign out[1172] = layer_0[1657] ^ layer_0[2285]; 
    assign out[1173] = layer_0[107] ^ layer_0[1645]; 
    assign out[1174] = ~(layer_0[1736] ^ layer_0[2063]); 
    assign out[1175] = layer_0[681] ^ layer_0[2160]; 
    assign out[1176] = layer_0[2044] | layer_0[2011]; 
    assign out[1177] = ~layer_0[829] | (layer_0[829] & layer_0[615]); 
    assign out[1178] = ~(layer_0[1179] ^ layer_0[497]); 
    assign out[1179] = layer_0[537] ^ layer_0[700]; 
    assign out[1180] = ~(layer_0[87] ^ layer_0[1194]); 
    assign out[1181] = ~layer_0[2349]; 
    assign out[1182] = layer_0[1114] ^ layer_0[1792]; 
    assign out[1183] = ~(layer_0[2102] | layer_0[1067]); 
    assign out[1184] = layer_0[2187] ^ layer_0[2472]; 
    assign out[1185] = layer_0[2502]; 
    assign out[1186] = ~(layer_0[821] ^ layer_0[949]); 
    assign out[1187] = layer_0[1698] & layer_0[383]; 
    assign out[1188] = layer_0[2416] ^ layer_0[1549]; 
    assign out[1189] = layer_0[589]; 
    assign out[1190] = ~layer_0[728]; 
    assign out[1191] = ~(layer_0[2444] | layer_0[1251]); 
    assign out[1192] = layer_0[1250]; 
    assign out[1193] = layer_0[2088] & ~layer_0[147]; 
    assign out[1194] = layer_0[705] | layer_0[2128]; 
    assign out[1195] = ~layer_0[2227]; 
    assign out[1196] = layer_0[47] & ~layer_0[1693]; 
    assign out[1197] = layer_0[2099] & ~layer_0[252]; 
    assign out[1198] = ~(layer_0[1535] ^ layer_0[346]); 
    assign out[1199] = layer_0[1337]; 
    assign out[1200] = layer_0[1644] | layer_0[1197]; 
    assign out[1201] = layer_0[2545] | layer_0[947]; 
    assign out[1202] = layer_0[1781] & ~layer_0[1926]; 
    assign out[1203] = layer_0[445] ^ layer_0[2069]; 
    assign out[1204] = layer_0[1368] & ~layer_0[960]; 
    assign out[1205] = layer_0[299] ^ layer_0[918]; 
    assign out[1206] = layer_0[2440] ^ layer_0[2174]; 
    assign out[1207] = ~(layer_0[525] ^ layer_0[1678]); 
    assign out[1208] = layer_0[1310] & layer_0[2151]; 
    assign out[1209] = ~layer_0[545]; 
    assign out[1210] = ~(layer_0[992] ^ layer_0[962]); 
    assign out[1211] = layer_0[2139] & ~layer_0[2343]; 
    assign out[1212] = ~(layer_0[2283] | layer_0[1232]); 
    assign out[1213] = layer_0[894] ^ layer_0[2159]; 
    assign out[1214] = layer_0[588] & layer_0[1639]; 
    assign out[1215] = layer_0[1560] ^ layer_0[776]; 
    assign out[1216] = layer_0[1004] ^ layer_0[79]; 
    assign out[1217] = layer_0[62] & layer_0[1687]; 
    assign out[1218] = layer_0[2542] & ~layer_0[1060]; 
    assign out[1219] = layer_0[1031] & ~layer_0[1581]; 
    assign out[1220] = layer_0[1352] ^ layer_0[495]; 
    assign out[1221] = layer_0[2257] ^ layer_0[336]; 
    assign out[1222] = ~(layer_0[1539] ^ layer_0[1005]); 
    assign out[1223] = layer_0[2242]; 
    assign out[1224] = ~(layer_0[1402] ^ layer_0[1286]); 
    assign out[1225] = layer_0[741] & ~layer_0[1734]; 
    assign out[1226] = layer_0[998] ^ layer_0[165]; 
    assign out[1227] = layer_0[2040] | layer_0[1263]; 
    assign out[1228] = ~(layer_0[230] ^ layer_0[2043]); 
    assign out[1229] = ~(layer_0[688] | layer_0[1971]); 
    assign out[1230] = layer_0[1246] & ~layer_0[221]; 
    assign out[1231] = ~(layer_0[530] ^ layer_0[2525]); 
    assign out[1232] = layer_0[730] & ~layer_0[1975]; 
    assign out[1233] = ~layer_0[1312]; 
    assign out[1234] = ~(layer_0[1024] | layer_0[653]); 
    assign out[1235] = ~(layer_0[68] & layer_0[401]); 
    assign out[1236] = layer_0[178] & ~layer_0[1335]; 
    assign out[1237] = layer_0[846] ^ layer_0[2056]; 
    assign out[1238] = layer_0[2104]; 
    assign out[1239] = ~layer_0[1347]; 
    assign out[1240] = layer_0[580] ^ layer_0[2025]; 
    assign out[1241] = ~(layer_0[1604] ^ layer_0[1671]); 
    assign out[1242] = ~(layer_0[832] ^ layer_0[1755]); 
    assign out[1243] = layer_0[1339] & ~layer_0[1715]; 
    assign out[1244] = ~(layer_0[1516] ^ layer_0[2392]); 
    assign out[1245] = layer_0[1424] | layer_0[2512]; 
    assign out[1246] = ~layer_0[915] | (layer_0[1764] & layer_0[915]); 
    assign out[1247] = layer_0[510] & layer_0[1426]; 
    assign out[1248] = layer_0[326] & layer_0[226]; 
    assign out[1249] = layer_0[899] & ~layer_0[478]; 
    assign out[1250] = ~(layer_0[711] ^ layer_0[1284]); 
    assign out[1251] = layer_0[908] ^ layer_0[1086]; 
    assign out[1252] = ~(layer_0[1590] ^ layer_0[602]); 
    assign out[1253] = ~layer_0[1441]; 
    assign out[1254] = ~layer_0[2315]; 
    assign out[1255] = ~layer_0[1328]; 
    assign out[1256] = layer_0[1948] ^ layer_0[1551]; 
    assign out[1257] = layer_0[1482]; 
    assign out[1258] = layer_0[750] & ~layer_0[2450]; 
    assign out[1259] = ~layer_0[716]; 
    assign out[1260] = ~(layer_0[932] ^ layer_0[797]); 
    assign out[1261] = layer_0[1936]; 
    assign out[1262] = layer_0[1999] ^ layer_0[569]; 
    assign out[1263] = layer_0[2442]; 
    assign out[1264] = layer_0[1600] ^ layer_0[283]; 
    assign out[1265] = ~layer_0[2402]; 
    assign out[1266] = layer_0[868]; 
    assign out[1267] = layer_0[2342] ^ layer_0[1178]; 
    assign out[1268] = layer_0[2550] & layer_0[1301]; 
    assign out[1269] = layer_0[1483] & ~layer_0[458]; 
    assign out[1270] = 1'b0; 
    assign out[1271] = 1'b0; 
    assign out[1272] = 1'b0; 
    assign out[1273] = 1'b0; 
    assign out[1274] = 1'b0; 
    assign out[1275] = 1'b0; 
    assign out[1276] = 1'b0; 
    assign out[1277] = 1'b0; 
    assign out[1278] = 1'b0; 
    assign out[1279] = 1'b0; 
    assign out[1280] = 1'b0; 
    assign out[1281] = 1'b0; 
    assign out[1282] = 1'b0; 
    assign out[1283] = 1'b0; 
    assign out[1284] = 1'b0; 
    assign out[1285] = 1'b0; 
    assign out[1286] = 1'b0; 
    assign out[1287] = 1'b0; 
    assign out[1288] = 1'b0; 
    assign out[1289] = 1'b0; 
    assign out[1290] = 1'b0; 
    assign out[1291] = 1'b0; 
    assign out[1292] = 1'b0; 
    assign out[1293] = 1'b0; 
    assign out[1294] = 1'b0; 
    assign out[1295] = 1'b0; 
    assign out[1296] = 1'b0; 
    assign out[1297] = 1'b0; 
    assign out[1298] = 1'b0; 
    assign out[1299] = 1'b0; 
    assign out[1300] = 1'b0; 
    assign out[1301] = 1'b0; 
    assign out[1302] = 1'b0; 
    assign out[1303] = 1'b0; 
    assign out[1304] = 1'b0; 
    assign out[1305] = 1'b0; 
    assign out[1306] = 1'b0; 
    assign out[1307] = 1'b0; 
    assign out[1308] = 1'b0; 
    assign out[1309] = 1'b0; 
    assign out[1310] = 1'b0; 
    assign out[1311] = 1'b0; 
    assign out[1312] = 1'b0; 
    assign out[1313] = 1'b0; 
    assign out[1314] = 1'b0; 
    assign out[1315] = 1'b0; 
    assign out[1316] = 1'b0; 
    assign out[1317] = 1'b0; 
    assign out[1318] = 1'b0; 
    assign out[1319] = 1'b0; 
    assign out[1320] = 1'b0; 
    assign out[1321] = 1'b0; 
    assign out[1322] = 1'b0; 
    assign out[1323] = 1'b0; 
    assign out[1324] = 1'b0; 
    assign out[1325] = 1'b0; 
    assign out[1326] = 1'b0; 
    assign out[1327] = 1'b0; 
    assign out[1328] = 1'b0; 
    assign out[1329] = 1'b0; 
    assign out[1330] = 1'b0; 
    assign out[1331] = 1'b0; 
    assign out[1332] = 1'b0; 
    assign out[1333] = 1'b0; 
    assign out[1334] = 1'b0; 
    assign out[1335] = 1'b0; 
    assign out[1336] = 1'b0; 
    assign out[1337] = 1'b0; 
    assign out[1338] = 1'b0; 
    assign out[1339] = 1'b0; 
    assign out[1340] = 1'b0; 
    assign out[1341] = 1'b0; 
    assign out[1342] = 1'b0; 
    assign out[1343] = 1'b0; 
    assign out[1344] = 1'b0; 
    assign out[1345] = 1'b0; 
    assign out[1346] = 1'b0; 
    assign out[1347] = 1'b0; 
    assign out[1348] = 1'b0; 
    assign out[1349] = 1'b0; 
    assign out[1350] = 1'b0; 
    assign out[1351] = 1'b0; 
    assign out[1352] = 1'b0; 
    assign out[1353] = 1'b0; 
    assign out[1354] = 1'b0; 
    assign out[1355] = 1'b0; 
    assign out[1356] = 1'b0; 
    assign out[1357] = 1'b0; 
    assign out[1358] = 1'b0; 
    assign out[1359] = 1'b0; 
    assign out[1360] = 1'b0; 
    assign out[1361] = 1'b0; 
    assign out[1362] = 1'b0; 
    assign out[1363] = 1'b0; 
    assign out[1364] = 1'b0; 
    assign out[1365] = 1'b0; 
    assign out[1366] = 1'b0; 
    assign out[1367] = 1'b0; 
    assign out[1368] = 1'b0; 
    assign out[1369] = 1'b0; 
    assign out[1370] = 1'b0; 
    assign out[1371] = 1'b0; 
    assign out[1372] = 1'b0; 
    assign out[1373] = 1'b0; 
    assign out[1374] = 1'b0; 
    assign out[1375] = 1'b0; 
    assign out[1376] = 1'b0; 
    assign out[1377] = 1'b0; 
    assign out[1378] = 1'b0; 
    assign out[1379] = 1'b0; 
    assign out[1380] = 1'b0; 
    assign out[1381] = 1'b0; 
    assign out[1382] = 1'b0; 
    assign out[1383] = 1'b0; 
    assign out[1384] = 1'b0; 
    assign out[1385] = 1'b0; 
    assign out[1386] = 1'b0; 
    assign out[1387] = 1'b0; 
    assign out[1388] = 1'b0; 
    assign out[1389] = 1'b0; 
    assign out[1390] = 1'b0; 
    assign out[1391] = 1'b0; 
    assign out[1392] = 1'b0; 
    assign out[1393] = 1'b0; 
    assign out[1394] = 1'b0; 
    assign out[1395] = 1'b0; 
    assign out[1396] = 1'b0; 
    assign out[1397] = 1'b0; 
    assign out[1398] = 1'b0; 
    assign out[1399] = 1'b0; 
    assign out[1400] = 1'b0; 
    assign out[1401] = 1'b0; 
    assign out[1402] = 1'b0; 
    assign out[1403] = 1'b0; 
    assign out[1404] = 1'b0; 
    assign out[1405] = 1'b0; 
    assign out[1406] = 1'b0; 
    assign out[1407] = 1'b0; 
    assign out[1408] = 1'b0; 
    assign out[1409] = 1'b0; 
    assign out[1410] = 1'b0; 
    assign out[1411] = 1'b0; 
    assign out[1412] = 1'b0; 
    assign out[1413] = 1'b0; 
    assign out[1414] = 1'b0; 
    assign out[1415] = 1'b0; 
    assign out[1416] = 1'b0; 
    assign out[1417] = 1'b0; 
    assign out[1418] = 1'b0; 
    assign out[1419] = 1'b0; 
    assign out[1420] = 1'b0; 
    assign out[1421] = 1'b0; 
    assign out[1422] = 1'b0; 
    assign out[1423] = 1'b0; 
    assign out[1424] = 1'b0; 
    assign out[1425] = 1'b0; 
    assign out[1426] = 1'b0; 
    assign out[1427] = 1'b0; 
    assign out[1428] = 1'b0; 
    assign out[1429] = 1'b0; 
    assign out[1430] = 1'b0; 
    assign out[1431] = 1'b0; 
    assign out[1432] = 1'b0; 
    assign out[1433] = 1'b0; 
    assign out[1434] = 1'b0; 
    assign out[1435] = 1'b0; 
    assign out[1436] = 1'b0; 
    assign out[1437] = 1'b0; 
    assign out[1438] = 1'b0; 
    assign out[1439] = 1'b0; 
    assign out[1440] = 1'b0; 
    assign out[1441] = 1'b0; 
    assign out[1442] = 1'b0; 
    assign out[1443] = 1'b0; 
    assign out[1444] = 1'b0; 
    assign out[1445] = 1'b0; 
    assign out[1446] = 1'b0; 
    assign out[1447] = 1'b0; 
    assign out[1448] = 1'b0; 
    assign out[1449] = 1'b0; 
    assign out[1450] = 1'b0; 
    assign out[1451] = 1'b0; 
    assign out[1452] = 1'b0; 
    assign out[1453] = 1'b0; 
    assign out[1454] = 1'b0; 
    assign out[1455] = 1'b0; 
    assign out[1456] = 1'b0; 
    assign out[1457] = 1'b0; 
    assign out[1458] = 1'b0; 
    assign out[1459] = 1'b0; 
    assign out[1460] = 1'b0; 
    assign out[1461] = 1'b0; 
    assign out[1462] = 1'b0; 
    assign out[1463] = 1'b0; 
    assign out[1464] = 1'b0; 
    assign out[1465] = 1'b0; 
    assign out[1466] = 1'b0; 
    assign out[1467] = 1'b0; 
    assign out[1468] = 1'b0; 
    assign out[1469] = 1'b0; 
    assign out[1470] = 1'b0; 
    assign out[1471] = 1'b0; 
    assign out[1472] = 1'b0; 
    assign out[1473] = 1'b0; 
    assign out[1474] = 1'b0; 
    assign out[1475] = 1'b0; 
    assign out[1476] = 1'b0; 
    assign out[1477] = 1'b0; 
    assign out[1478] = 1'b0; 
    assign out[1479] = 1'b0; 
    assign out[1480] = 1'b0; 
    assign out[1481] = 1'b0; 
    assign out[1482] = 1'b0; 
    assign out[1483] = 1'b0; 
    assign out[1484] = 1'b0; 
    assign out[1485] = 1'b0; 
    assign out[1486] = 1'b0; 
    assign out[1487] = 1'b0; 
    assign out[1488] = 1'b0; 
    assign out[1489] = 1'b0; 
    assign out[1490] = 1'b0; 
    assign out[1491] = 1'b0; 
    assign out[1492] = 1'b0; 
    assign out[1493] = 1'b0; 
    assign out[1494] = 1'b0; 
    assign out[1495] = 1'b0; 
    assign out[1496] = 1'b0; 
    assign out[1497] = 1'b0; 
    assign out[1498] = 1'b0; 
    assign out[1499] = 1'b0; 
    assign out[1500] = 1'b0; 
    assign out[1501] = 1'b0; 
    assign out[1502] = 1'b0; 
    assign out[1503] = 1'b0; 
    assign out[1504] = 1'b0; 
    assign out[1505] = 1'b0; 
    assign out[1506] = 1'b0; 
    assign out[1507] = 1'b0; 
    assign out[1508] = 1'b0; 
    assign out[1509] = 1'b0; 
    assign out[1510] = 1'b0; 
    assign out[1511] = 1'b0; 
    assign out[1512] = 1'b0; 
    assign out[1513] = 1'b0; 
    assign out[1514] = 1'b0; 
    assign out[1515] = 1'b0; 
    assign out[1516] = 1'b0; 
    assign out[1517] = 1'b0; 
    assign out[1518] = 1'b0; 
    assign out[1519] = 1'b0; 
    assign out[1520] = 1'b0; 
    assign out[1521] = 1'b0; 
    assign out[1522] = 1'b0; 
    assign out[1523] = 1'b0; 
    assign out[1524] = 1'b0; 
    assign out[1525] = 1'b0; 
    assign out[1526] = 1'b0; 
    assign out[1527] = 1'b0; 
    assign out[1528] = 1'b0; 
    assign out[1529] = 1'b0; 
    assign out[1530] = 1'b0; 
    assign out[1531] = 1'b0; 
    assign out[1532] = 1'b0; 
    assign out[1533] = 1'b0; 
    assign out[1534] = 1'b0; 
    assign out[1535] = 1'b0; 
    assign out[1536] = 1'b0; 
    assign out[1537] = 1'b0; 
    assign out[1538] = 1'b0; 
    assign out[1539] = 1'b0; 
    assign out[1540] = 1'b0; 
    assign out[1541] = 1'b0; 
    assign out[1542] = 1'b0; 
    assign out[1543] = 1'b0; 
    assign out[1544] = 1'b0; 
    assign out[1545] = 1'b0; 
    assign out[1546] = 1'b0; 
    assign out[1547] = 1'b0; 
    assign out[1548] = 1'b0; 
    assign out[1549] = 1'b0; 
    assign out[1550] = 1'b0; 
    assign out[1551] = 1'b0; 
    assign out[1552] = 1'b0; 
    assign out[1553] = 1'b0; 
    assign out[1554] = 1'b0; 
    assign out[1555] = 1'b0; 
    assign out[1556] = 1'b0; 
    assign out[1557] = 1'b0; 
    assign out[1558] = 1'b0; 
    assign out[1559] = 1'b0; 
    assign out[1560] = 1'b0; 
    assign out[1561] = 1'b0; 
    assign out[1562] = 1'b0; 
    assign out[1563] = 1'b0; 
    assign out[1564] = 1'b0; 
    assign out[1565] = 1'b0; 
    assign out[1566] = 1'b0; 
    assign out[1567] = 1'b0; 
    assign out[1568] = 1'b0; 
    assign out[1569] = 1'b0; 
    assign out[1570] = 1'b0; 
    assign out[1571] = 1'b0; 
    assign out[1572] = 1'b0; 
    assign out[1573] = 1'b0; 
    assign out[1574] = 1'b0; 
    assign out[1575] = 1'b0; 
    assign out[1576] = 1'b0; 
    assign out[1577] = 1'b0; 
    assign out[1578] = 1'b0; 
    assign out[1579] = 1'b0; 
    assign out[1580] = 1'b0; 
    assign out[1581] = 1'b0; 
    assign out[1582] = 1'b0; 
    assign out[1583] = 1'b0; 
    assign out[1584] = 1'b0; 
    assign out[1585] = 1'b0; 
    assign out[1586] = 1'b0; 
    assign out[1587] = 1'b0; 
    assign out[1588] = 1'b0; 
    assign out[1589] = 1'b0; 
    assign out[1590] = 1'b0; 
    assign out[1591] = 1'b0; 
    assign out[1592] = 1'b0; 
    assign out[1593] = 1'b0; 
    assign out[1594] = 1'b0; 
    assign out[1595] = 1'b0; 
    assign out[1596] = 1'b0; 
    assign out[1597] = 1'b0; 
    assign out[1598] = 1'b0; 
    assign out[1599] = 1'b0; 
    assign out[1600] = 1'b0; 
    assign out[1601] = 1'b0; 
    assign out[1602] = 1'b0; 
    assign out[1603] = 1'b0; 
    assign out[1604] = 1'b0; 
    assign out[1605] = 1'b0; 
    assign out[1606] = 1'b0; 
    assign out[1607] = 1'b0; 
    assign out[1608] = 1'b0; 
    assign out[1609] = 1'b0; 
    assign out[1610] = 1'b0; 
    assign out[1611] = 1'b0; 
    assign out[1612] = 1'b0; 
    assign out[1613] = 1'b0; 
    assign out[1614] = 1'b0; 
    assign out[1615] = 1'b0; 
    assign out[1616] = 1'b0; 
    assign out[1617] = 1'b0; 
    assign out[1618] = 1'b0; 
    assign out[1619] = 1'b0; 
    assign out[1620] = 1'b0; 
    assign out[1621] = 1'b0; 
    assign out[1622] = 1'b0; 
    assign out[1623] = 1'b0; 
    assign out[1624] = 1'b0; 
    assign out[1625] = 1'b0; 
    assign out[1626] = 1'b0; 
    assign out[1627] = 1'b0; 
    assign out[1628] = 1'b0; 
    assign out[1629] = 1'b0; 
    assign out[1630] = 1'b0; 
    assign out[1631] = 1'b0; 
    assign out[1632] = 1'b0; 
    assign out[1633] = 1'b0; 
    assign out[1634] = 1'b0; 
    assign out[1635] = 1'b0; 
    assign out[1636] = 1'b0; 
    assign out[1637] = 1'b0; 
    assign out[1638] = 1'b0; 
    assign out[1639] = 1'b0; 
    assign out[1640] = 1'b0; 
    assign out[1641] = 1'b0; 
    assign out[1642] = 1'b0; 
    assign out[1643] = 1'b0; 
    assign out[1644] = 1'b0; 
    assign out[1645] = 1'b0; 
    assign out[1646] = 1'b0; 
    assign out[1647] = 1'b0; 
    assign out[1648] = 1'b0; 
    assign out[1649] = 1'b0; 
    assign out[1650] = 1'b0; 
    assign out[1651] = 1'b0; 
    assign out[1652] = 1'b0; 
    assign out[1653] = 1'b0; 
    assign out[1654] = 1'b0; 
    assign out[1655] = 1'b0; 
    assign out[1656] = 1'b0; 
    assign out[1657] = 1'b0; 
    assign out[1658] = 1'b0; 
    assign out[1659] = 1'b0; 
    assign out[1660] = 1'b0; 
    assign out[1661] = 1'b0; 
    assign out[1662] = 1'b0; 
    assign out[1663] = 1'b0; 
    assign out[1664] = 1'b0; 
    assign out[1665] = 1'b0; 
    assign out[1666] = 1'b0; 
    assign out[1667] = 1'b0; 
    assign out[1668] = 1'b0; 
    assign out[1669] = 1'b0; 
    assign out[1670] = 1'b0; 
    assign out[1671] = 1'b0; 
    assign out[1672] = 1'b0; 
    assign out[1673] = 1'b0; 
    assign out[1674] = 1'b0; 
    assign out[1675] = 1'b0; 
    assign out[1676] = 1'b0; 
    assign out[1677] = 1'b0; 
    assign out[1678] = 1'b0; 
    assign out[1679] = 1'b0; 
    assign out[1680] = 1'b0; 
    assign out[1681] = 1'b0; 
    assign out[1682] = 1'b0; 
    assign out[1683] = 1'b0; 
    assign out[1684] = 1'b0; 
    assign out[1685] = 1'b0; 
    assign out[1686] = 1'b0; 
    assign out[1687] = 1'b0; 
    assign out[1688] = 1'b0; 
    assign out[1689] = 1'b0; 
    assign out[1690] = 1'b0; 
    assign out[1691] = 1'b0; 
    assign out[1692] = 1'b0; 
    assign out[1693] = 1'b0; 
    assign out[1694] = 1'b0; 
    assign out[1695] = 1'b0; 
    assign out[1696] = 1'b0; 
    assign out[1697] = 1'b0; 
    assign out[1698] = 1'b0; 
    assign out[1699] = 1'b0; 
    assign out[1700] = 1'b0; 
    assign out[1701] = 1'b0; 
    assign out[1702] = 1'b0; 
    assign out[1703] = 1'b0; 
    assign out[1704] = 1'b0; 
    assign out[1705] = 1'b0; 
    assign out[1706] = 1'b0; 
    assign out[1707] = 1'b0; 
    assign out[1708] = 1'b0; 
    assign out[1709] = 1'b0; 
    assign out[1710] = 1'b0; 
    assign out[1711] = 1'b0; 
    assign out[1712] = 1'b0; 
    assign out[1713] = 1'b0; 
    assign out[1714] = 1'b0; 
    assign out[1715] = 1'b0; 
    assign out[1716] = 1'b0; 
    assign out[1717] = 1'b0; 
    assign out[1718] = 1'b0; 
    assign out[1719] = 1'b0; 
    assign out[1720] = 1'b0; 
    assign out[1721] = 1'b0; 
    assign out[1722] = 1'b0; 
    assign out[1723] = 1'b0; 
    assign out[1724] = 1'b0; 
    assign out[1725] = 1'b0; 
    assign out[1726] = 1'b0; 
    assign out[1727] = 1'b0; 
    assign out[1728] = 1'b0; 
    assign out[1729] = 1'b0; 
    assign out[1730] = 1'b0; 
    assign out[1731] = 1'b0; 
    assign out[1732] = 1'b0; 
    assign out[1733] = 1'b0; 
    assign out[1734] = 1'b0; 
    assign out[1735] = 1'b0; 
    assign out[1736] = 1'b0; 
    assign out[1737] = 1'b0; 
    assign out[1738] = 1'b0; 
    assign out[1739] = 1'b0; 
    assign out[1740] = 1'b0; 
    assign out[1741] = 1'b0; 
    assign out[1742] = 1'b0; 
    assign out[1743] = 1'b0; 
    assign out[1744] = 1'b0; 
    assign out[1745] = 1'b0; 
    assign out[1746] = 1'b0; 
    assign out[1747] = 1'b0; 
    assign out[1748] = 1'b0; 
    assign out[1749] = 1'b0; 
    assign out[1750] = 1'b0; 
    assign out[1751] = 1'b0; 
    assign out[1752] = 1'b0; 
    assign out[1753] = 1'b0; 
    assign out[1754] = 1'b0; 
    assign out[1755] = 1'b0; 
    assign out[1756] = 1'b0; 
    assign out[1757] = 1'b0; 
    assign out[1758] = 1'b0; 
    assign out[1759] = 1'b0; 
    assign out[1760] = 1'b0; 
    assign out[1761] = 1'b0; 
    assign out[1762] = 1'b0; 
    assign out[1763] = 1'b0; 
    assign out[1764] = 1'b0; 
    assign out[1765] = 1'b0; 
    assign out[1766] = 1'b0; 
    assign out[1767] = 1'b0; 
    assign out[1768] = 1'b0; 
    assign out[1769] = 1'b0; 
    assign out[1770] = 1'b0; 
    assign out[1771] = 1'b0; 
    assign out[1772] = 1'b0; 
    assign out[1773] = 1'b0; 
    assign out[1774] = 1'b0; 
    assign out[1775] = 1'b0; 
    assign out[1776] = 1'b0; 
    assign out[1777] = 1'b0; 
    assign out[1778] = 1'b0; 
    assign out[1779] = 1'b0; 
    assign out[1780] = 1'b0; 
    assign out[1781] = 1'b0; 
    assign out[1782] = 1'b0; 
    assign out[1783] = 1'b0; 
    assign out[1784] = 1'b0; 
    assign out[1785] = 1'b0; 
    assign out[1786] = 1'b0; 
    assign out[1787] = 1'b0; 
    assign out[1788] = 1'b0; 
    assign out[1789] = 1'b0; 
    assign out[1790] = 1'b0; 
    assign out[1791] = 1'b0; 
    assign out[1792] = 1'b0; 
    assign out[1793] = 1'b0; 
    assign out[1794] = 1'b0; 
    assign out[1795] = 1'b0; 
    assign out[1796] = 1'b0; 
    assign out[1797] = 1'b0; 
    assign out[1798] = 1'b0; 
    assign out[1799] = 1'b0; 
    assign out[1800] = 1'b0; 
    assign out[1801] = 1'b0; 
    assign out[1802] = 1'b0; 
    assign out[1803] = 1'b0; 
    assign out[1804] = 1'b0; 
    assign out[1805] = 1'b0; 
    assign out[1806] = 1'b0; 
    assign out[1807] = 1'b0; 
    assign out[1808] = 1'b0; 
    assign out[1809] = 1'b0; 
    assign out[1810] = 1'b0; 
    assign out[1811] = 1'b0; 
    assign out[1812] = 1'b0; 
    assign out[1813] = 1'b0; 
    assign out[1814] = 1'b0; 
    assign out[1815] = 1'b0; 
    assign out[1816] = 1'b0; 
    assign out[1817] = 1'b0; 
    assign out[1818] = 1'b0; 
    assign out[1819] = 1'b0; 
    assign out[1820] = 1'b0; 
    assign out[1821] = 1'b0; 
    assign out[1822] = 1'b0; 
    assign out[1823] = 1'b0; 
    assign out[1824] = 1'b0; 
    assign out[1825] = 1'b0; 
    assign out[1826] = 1'b0; 
    assign out[1827] = 1'b0; 
    assign out[1828] = 1'b0; 
    assign out[1829] = 1'b0; 
    assign out[1830] = 1'b0; 
    assign out[1831] = 1'b0; 
    assign out[1832] = 1'b0; 
    assign out[1833] = 1'b0; 
    assign out[1834] = 1'b0; 
    assign out[1835] = 1'b0; 
    assign out[1836] = 1'b0; 
    assign out[1837] = 1'b0; 
    assign out[1838] = 1'b0; 
    assign out[1839] = 1'b0; 
    assign out[1840] = 1'b0; 
    assign out[1841] = 1'b0; 
    assign out[1842] = 1'b0; 
    assign out[1843] = 1'b0; 
    assign out[1844] = 1'b0; 
    assign out[1845] = 1'b0; 
    assign out[1846] = 1'b0; 
    assign out[1847] = 1'b0; 
    assign out[1848] = 1'b0; 
    assign out[1849] = 1'b0; 
    assign out[1850] = 1'b0; 
    assign out[1851] = 1'b0; 
    assign out[1852] = 1'b0; 
    assign out[1853] = 1'b0; 
    assign out[1854] = 1'b0; 
    assign out[1855] = 1'b0; 
    assign out[1856] = 1'b0; 
    assign out[1857] = 1'b0; 
    assign out[1858] = 1'b0; 
    assign out[1859] = 1'b0; 
    assign out[1860] = 1'b0; 
    assign out[1861] = 1'b0; 
    assign out[1862] = 1'b0; 
    assign out[1863] = 1'b0; 
    assign out[1864] = 1'b0; 
    assign out[1865] = 1'b0; 
    assign out[1866] = 1'b0; 
    assign out[1867] = 1'b0; 
    assign out[1868] = 1'b0; 
    assign out[1869] = 1'b0; 
    assign out[1870] = 1'b0; 
    assign out[1871] = 1'b0; 
    assign out[1872] = 1'b0; 
    assign out[1873] = 1'b0; 
    assign out[1874] = 1'b0; 
    assign out[1875] = 1'b0; 
    assign out[1876] = 1'b0; 
    assign out[1877] = 1'b0; 
    assign out[1878] = 1'b0; 
    assign out[1879] = 1'b0; 
    assign out[1880] = 1'b0; 
    assign out[1881] = 1'b0; 
    assign out[1882] = 1'b0; 
    assign out[1883] = 1'b0; 
    assign out[1884] = 1'b0; 
    assign out[1885] = 1'b0; 
    assign out[1886] = 1'b0; 
    assign out[1887] = 1'b0; 
    assign out[1888] = 1'b0; 
    assign out[1889] = 1'b0; 
    assign out[1890] = 1'b0; 
    assign out[1891] = 1'b0; 
    assign out[1892] = 1'b0; 
    assign out[1893] = 1'b0; 
    assign out[1894] = 1'b0; 
    assign out[1895] = 1'b0; 
    assign out[1896] = 1'b0; 
    assign out[1897] = 1'b0; 
    assign out[1898] = 1'b0; 
    assign out[1899] = 1'b0; 
    assign out[1900] = 1'b0; 
    assign out[1901] = 1'b0; 
    assign out[1902] = 1'b0; 
    assign out[1903] = 1'b0; 
    assign out[1904] = 1'b0; 
    assign out[1905] = 1'b0; 
    assign out[1906] = 1'b0; 
    assign out[1907] = 1'b0; 
    assign out[1908] = 1'b0; 
    assign out[1909] = 1'b0; 
    assign out[1910] = 1'b0; 
    assign out[1911] = 1'b0; 
    assign out[1912] = 1'b0; 
    assign out[1913] = 1'b0; 
    assign out[1914] = 1'b0; 
    assign out[1915] = 1'b0; 
    assign out[1916] = 1'b0; 
    assign out[1917] = 1'b0; 
    assign out[1918] = 1'b0; 
    assign out[1919] = 1'b0; 
    assign out[1920] = 1'b0; 
    assign out[1921] = 1'b0; 
    assign out[1922] = 1'b0; 
    assign out[1923] = 1'b0; 
    assign out[1924] = 1'b0; 
    assign out[1925] = 1'b0; 
    assign out[1926] = 1'b0; 
    assign out[1927] = 1'b0; 
    assign out[1928] = 1'b0; 
    assign out[1929] = 1'b0; 
    assign out[1930] = 1'b0; 
    assign out[1931] = 1'b0; 
    assign out[1932] = 1'b0; 
    assign out[1933] = 1'b0; 
    assign out[1934] = 1'b0; 
    assign out[1935] = 1'b0; 
    assign out[1936] = 1'b0; 
    assign out[1937] = 1'b0; 
    assign out[1938] = 1'b0; 
    assign out[1939] = 1'b0; 
    assign out[1940] = 1'b0; 
    assign out[1941] = 1'b0; 
    assign out[1942] = 1'b0; 
    assign out[1943] = 1'b0; 
    assign out[1944] = 1'b0; 
    assign out[1945] = 1'b0; 
    assign out[1946] = 1'b0; 
    assign out[1947] = 1'b0; 
    assign out[1948] = 1'b0; 
    assign out[1949] = 1'b0; 
    assign out[1950] = 1'b0; 
    assign out[1951] = 1'b0; 
    assign out[1952] = 1'b0; 
    assign out[1953] = 1'b0; 
    assign out[1954] = 1'b0; 
    assign out[1955] = 1'b0; 
    assign out[1956] = 1'b0; 
    assign out[1957] = 1'b0; 
    assign out[1958] = 1'b0; 
    assign out[1959] = 1'b0; 
    assign out[1960] = 1'b0; 
    assign out[1961] = 1'b0; 
    assign out[1962] = 1'b0; 
    assign out[1963] = 1'b0; 
    assign out[1964] = 1'b0; 
    assign out[1965] = 1'b0; 
    assign out[1966] = 1'b0; 
    assign out[1967] = 1'b0; 
    assign out[1968] = 1'b0; 
    assign out[1969] = 1'b0; 
    assign out[1970] = 1'b0; 
    assign out[1971] = 1'b0; 
    assign out[1972] = 1'b0; 
    assign out[1973] = 1'b0; 
    assign out[1974] = 1'b0; 
    assign out[1975] = 1'b0; 
    assign out[1976] = 1'b0; 
    assign out[1977] = 1'b0; 
    assign out[1978] = 1'b0; 
    assign out[1979] = 1'b0; 
    assign out[1980] = 1'b0; 
    assign out[1981] = 1'b0; 
    assign out[1982] = 1'b0; 
    assign out[1983] = 1'b0; 
    assign out[1984] = 1'b0; 
    assign out[1985] = 1'b0; 
    assign out[1986] = 1'b0; 
    assign out[1987] = 1'b0; 
    assign out[1988] = 1'b0; 
    assign out[1989] = 1'b0; 
    assign out[1990] = 1'b0; 
    assign out[1991] = 1'b0; 
    assign out[1992] = 1'b0; 
    assign out[1993] = 1'b0; 
    assign out[1994] = 1'b0; 
    assign out[1995] = 1'b0; 
    assign out[1996] = 1'b0; 
    assign out[1997] = 1'b0; 
    assign out[1998] = 1'b0; 
    assign out[1999] = 1'b0; 
    assign out[2000] = 1'b0; 
    assign out[2001] = 1'b0; 
    assign out[2002] = 1'b0; 
    assign out[2003] = 1'b0; 
    assign out[2004] = 1'b0; 
    assign out[2005] = 1'b0; 
    assign out[2006] = 1'b0; 
    assign out[2007] = 1'b0; 
    assign out[2008] = 1'b0; 
    assign out[2009] = 1'b0; 
    assign out[2010] = 1'b0; 
    assign out[2011] = 1'b0; 
    assign out[2012] = 1'b0; 
    assign out[2013] = 1'b0; 
    assign out[2014] = 1'b0; 
    assign out[2015] = 1'b0; 
    assign out[2016] = 1'b0; 
    assign out[2017] = 1'b0; 
    assign out[2018] = 1'b0; 
    assign out[2019] = 1'b0; 
    assign out[2020] = 1'b0; 
    assign out[2021] = 1'b0; 
    assign out[2022] = 1'b0; 
    assign out[2023] = 1'b0; 
    assign out[2024] = 1'b0; 
    assign out[2025] = 1'b0; 
    assign out[2026] = 1'b0; 
    assign out[2027] = 1'b0; 
    assign out[2028] = 1'b0; 
    assign out[2029] = 1'b0; 
    assign out[2030] = 1'b0; 
    assign out[2031] = 1'b0; 
    assign out[2032] = 1'b0; 
    assign out[2033] = 1'b0; 
    assign out[2034] = 1'b0; 
    assign out[2035] = 1'b0; 
    assign out[2036] = 1'b0; 
    assign out[2037] = 1'b0; 
    assign out[2038] = 1'b0; 
    assign out[2039] = 1'b0; 
    assign out[2040] = 1'b0; 
    assign out[2041] = 1'b0; 
    assign out[2042] = 1'b0; 
    assign out[2043] = 1'b0; 
    assign out[2044] = 1'b0; 
    assign out[2045] = 1'b0; 
    assign out[2046] = 1'b0; 
    assign out[2047] = 1'b0; 
    assign out[2048] = 1'b0; 
    assign out[2049] = 1'b0; 
    assign out[2050] = 1'b0; 
    assign out[2051] = 1'b0; 
    assign out[2052] = 1'b0; 
    assign out[2053] = 1'b0; 
    assign out[2054] = 1'b0; 
    assign out[2055] = 1'b0; 
    assign out[2056] = 1'b0; 
    assign out[2057] = 1'b0; 
    assign out[2058] = 1'b0; 
    assign out[2059] = 1'b0; 
    assign out[2060] = 1'b0; 
    assign out[2061] = 1'b0; 
    assign out[2062] = 1'b0; 
    assign out[2063] = 1'b0; 
    assign out[2064] = 1'b0; 
    assign out[2065] = 1'b0; 
    assign out[2066] = 1'b0; 
    assign out[2067] = 1'b0; 
    assign out[2068] = 1'b0; 
    assign out[2069] = 1'b0; 
    assign out[2070] = 1'b0; 
    assign out[2071] = 1'b0; 
    assign out[2072] = 1'b0; 
    assign out[2073] = 1'b0; 
    assign out[2074] = 1'b0; 
    assign out[2075] = 1'b0; 
    assign out[2076] = 1'b0; 
    assign out[2077] = 1'b0; 
    assign out[2078] = 1'b0; 
    assign out[2079] = 1'b0; 
    assign out[2080] = 1'b0; 
    assign out[2081] = 1'b0; 
    assign out[2082] = 1'b0; 
    assign out[2083] = 1'b0; 
    assign out[2084] = 1'b0; 
    assign out[2085] = 1'b0; 
    assign out[2086] = 1'b0; 
    assign out[2087] = 1'b0; 
    assign out[2088] = 1'b0; 
    assign out[2089] = 1'b0; 
    assign out[2090] = 1'b0; 
    assign out[2091] = 1'b0; 
    assign out[2092] = 1'b0; 
    assign out[2093] = 1'b0; 
    assign out[2094] = 1'b0; 
    assign out[2095] = 1'b0; 
    assign out[2096] = 1'b0; 
    assign out[2097] = 1'b0; 
    assign out[2098] = 1'b0; 
    assign out[2099] = 1'b0; 
    assign out[2100] = 1'b0; 
    assign out[2101] = 1'b0; 
    assign out[2102] = 1'b0; 
    assign out[2103] = 1'b0; 
    assign out[2104] = 1'b0; 
    assign out[2105] = 1'b0; 
    assign out[2106] = 1'b0; 
    assign out[2107] = 1'b0; 
    assign out[2108] = 1'b0; 
    assign out[2109] = 1'b0; 
    assign out[2110] = 1'b0; 
    assign out[2111] = 1'b0; 
    assign out[2112] = 1'b0; 
    assign out[2113] = 1'b0; 
    assign out[2114] = 1'b0; 
    assign out[2115] = 1'b0; 
    assign out[2116] = 1'b0; 
    assign out[2117] = 1'b0; 
    assign out[2118] = 1'b0; 
    assign out[2119] = 1'b0; 
    assign out[2120] = 1'b0; 
    assign out[2121] = 1'b0; 
    assign out[2122] = 1'b0; 
    assign out[2123] = 1'b0; 
    assign out[2124] = 1'b0; 
    assign out[2125] = 1'b0; 
    assign out[2126] = 1'b0; 
    assign out[2127] = 1'b0; 
    assign out[2128] = 1'b0; 
    assign out[2129] = 1'b0; 
    assign out[2130] = 1'b0; 
    assign out[2131] = 1'b0; 
    assign out[2132] = 1'b0; 
    assign out[2133] = 1'b0; 
    assign out[2134] = 1'b0; 
    assign out[2135] = 1'b0; 
    assign out[2136] = 1'b0; 
    assign out[2137] = 1'b0; 
    assign out[2138] = 1'b0; 
    assign out[2139] = 1'b0; 
    assign out[2140] = 1'b0; 
    assign out[2141] = 1'b0; 
    assign out[2142] = 1'b0; 
    assign out[2143] = 1'b0; 
    assign out[2144] = 1'b0; 
    assign out[2145] = 1'b0; 
    assign out[2146] = 1'b0; 
    assign out[2147] = 1'b0; 
    assign out[2148] = 1'b0; 
    assign out[2149] = 1'b0; 
    assign out[2150] = 1'b0; 
    assign out[2151] = 1'b0; 
    assign out[2152] = 1'b0; 
    assign out[2153] = 1'b0; 
    assign out[2154] = 1'b0; 
    assign out[2155] = 1'b0; 
    assign out[2156] = 1'b0; 
    assign out[2157] = 1'b0; 
    assign out[2158] = 1'b0; 
    assign out[2159] = 1'b0; 
    assign out[2160] = 1'b0; 
    assign out[2161] = 1'b0; 
    assign out[2162] = 1'b0; 
    assign out[2163] = 1'b0; 
    assign out[2164] = 1'b0; 
    assign out[2165] = 1'b0; 
    assign out[2166] = 1'b0; 
    assign out[2167] = 1'b0; 
    assign out[2168] = 1'b0; 
    assign out[2169] = 1'b0; 
    assign out[2170] = 1'b0; 
    assign out[2171] = 1'b0; 
    assign out[2172] = 1'b0; 
    assign out[2173] = 1'b0; 
    assign out[2174] = 1'b0; 
    assign out[2175] = 1'b0; 
    assign out[2176] = 1'b0; 
    assign out[2177] = 1'b0; 
    assign out[2178] = 1'b0; 
    assign out[2179] = 1'b0; 
    assign out[2180] = 1'b0; 
    assign out[2181] = 1'b0; 
    assign out[2182] = 1'b0; 
    assign out[2183] = 1'b0; 
    assign out[2184] = 1'b0; 
    assign out[2185] = 1'b0; 
    assign out[2186] = 1'b0; 
    assign out[2187] = 1'b0; 
    assign out[2188] = 1'b0; 
    assign out[2189] = 1'b0; 
    assign out[2190] = 1'b0; 
    assign out[2191] = 1'b0; 
    assign out[2192] = 1'b0; 
    assign out[2193] = 1'b0; 
    assign out[2194] = 1'b0; 
    assign out[2195] = 1'b0; 
    assign out[2196] = 1'b0; 
    assign out[2197] = 1'b0; 
    assign out[2198] = 1'b0; 
    assign out[2199] = 1'b0; 
    assign out[2200] = 1'b0; 
    assign out[2201] = 1'b0; 
    assign out[2202] = 1'b0; 
    assign out[2203] = 1'b0; 
    assign out[2204] = 1'b0; 
    assign out[2205] = 1'b0; 
    assign out[2206] = 1'b0; 
    assign out[2207] = 1'b0; 
    assign out[2208] = 1'b0; 
    assign out[2209] = 1'b0; 
    assign out[2210] = 1'b0; 
    assign out[2211] = 1'b0; 
    assign out[2212] = 1'b0; 
    assign out[2213] = 1'b0; 
    assign out[2214] = 1'b0; 
    assign out[2215] = 1'b0; 
    assign out[2216] = 1'b0; 
    assign out[2217] = 1'b0; 
    assign out[2218] = 1'b0; 
    assign out[2219] = 1'b0; 
    assign out[2220] = 1'b0; 
    assign out[2221] = 1'b0; 
    assign out[2222] = 1'b0; 
    assign out[2223] = 1'b0; 
    assign out[2224] = 1'b0; 
    assign out[2225] = 1'b0; 
    assign out[2226] = 1'b0; 
    assign out[2227] = 1'b0; 
    assign out[2228] = 1'b0; 
    assign out[2229] = 1'b0; 
    assign out[2230] = 1'b0; 
    assign out[2231] = 1'b0; 
    assign out[2232] = 1'b0; 
    assign out[2233] = 1'b0; 
    assign out[2234] = 1'b0; 
    assign out[2235] = 1'b0; 
    assign out[2236] = 1'b0; 
    assign out[2237] = 1'b0; 
    assign out[2238] = 1'b0; 
    assign out[2239] = 1'b0; 
    assign out[2240] = 1'b0; 
    assign out[2241] = 1'b0; 
    assign out[2242] = 1'b0; 
    assign out[2243] = 1'b0; 
    assign out[2244] = 1'b0; 
    assign out[2245] = 1'b0; 
    assign out[2246] = 1'b0; 
    assign out[2247] = 1'b0; 
    assign out[2248] = 1'b0; 
    assign out[2249] = 1'b0; 
    assign out[2250] = 1'b0; 
    assign out[2251] = 1'b0; 
    assign out[2252] = 1'b0; 
    assign out[2253] = 1'b0; 
    assign out[2254] = 1'b0; 
    assign out[2255] = 1'b0; 
    assign out[2256] = 1'b0; 
    assign out[2257] = 1'b0; 
    assign out[2258] = 1'b0; 
    assign out[2259] = 1'b0; 
    assign out[2260] = 1'b0; 
    assign out[2261] = 1'b0; 
    assign out[2262] = 1'b0; 
    assign out[2263] = 1'b0; 
    assign out[2264] = 1'b0; 
    assign out[2265] = 1'b0; 
    assign out[2266] = 1'b0; 
    assign out[2267] = 1'b0; 
    assign out[2268] = 1'b0; 
    assign out[2269] = 1'b0; 
    assign out[2270] = 1'b0; 
    assign out[2271] = 1'b0; 
    assign out[2272] = 1'b0; 
    assign out[2273] = 1'b0; 
    assign out[2274] = 1'b0; 
    assign out[2275] = 1'b0; 
    assign out[2276] = 1'b0; 
    assign out[2277] = 1'b0; 
    assign out[2278] = 1'b0; 
    assign out[2279] = 1'b0; 
    assign out[2280] = 1'b0; 
    assign out[2281] = 1'b0; 
    assign out[2282] = 1'b0; 
    assign out[2283] = 1'b0; 
    assign out[2284] = 1'b0; 
    assign out[2285] = 1'b0; 
    assign out[2286] = 1'b0; 
    assign out[2287] = 1'b0; 
    assign out[2288] = 1'b0; 
    assign out[2289] = 1'b0; 
    assign out[2290] = 1'b0; 
    assign out[2291] = 1'b0; 
    assign out[2292] = 1'b0; 
    assign out[2293] = 1'b0; 
    assign out[2294] = 1'b0; 
    assign out[2295] = 1'b0; 
    assign out[2296] = 1'b0; 
    assign out[2297] = 1'b0; 
    assign out[2298] = 1'b0; 
    assign out[2299] = 1'b0; 
    assign out[2300] = 1'b0; 
    assign out[2301] = 1'b0; 
    assign out[2302] = 1'b0; 
    assign out[2303] = 1'b0; 
    assign out[2304] = 1'b0; 
    assign out[2305] = 1'b0; 
    assign out[2306] = 1'b0; 
    assign out[2307] = 1'b0; 
    assign out[2308] = 1'b0; 
    assign out[2309] = 1'b0; 
    assign out[2310] = 1'b0; 
    assign out[2311] = 1'b0; 
    assign out[2312] = 1'b0; 
    assign out[2313] = 1'b0; 
    assign out[2314] = 1'b0; 
    assign out[2315] = 1'b0; 
    assign out[2316] = 1'b0; 
    assign out[2317] = 1'b0; 
    assign out[2318] = 1'b0; 
    assign out[2319] = 1'b0; 
    assign out[2320] = 1'b0; 
    assign out[2321] = 1'b0; 
    assign out[2322] = 1'b0; 
    assign out[2323] = 1'b0; 
    assign out[2324] = 1'b0; 
    assign out[2325] = 1'b0; 
    assign out[2326] = 1'b0; 
    assign out[2327] = 1'b0; 
    assign out[2328] = 1'b0; 
    assign out[2329] = 1'b0; 
    assign out[2330] = 1'b0; 
    assign out[2331] = 1'b0; 
    assign out[2332] = 1'b0; 
    assign out[2333] = 1'b0; 
    assign out[2334] = 1'b0; 
    assign out[2335] = 1'b0; 
    assign out[2336] = 1'b0; 
    assign out[2337] = 1'b0; 
    assign out[2338] = 1'b0; 
    assign out[2339] = 1'b0; 
    assign out[2340] = 1'b0; 
    assign out[2341] = 1'b0; 
    assign out[2342] = 1'b0; 
    assign out[2343] = 1'b0; 
    assign out[2344] = 1'b0; 
    assign out[2345] = 1'b0; 
    assign out[2346] = 1'b0; 
    assign out[2347] = 1'b0; 
    assign out[2348] = 1'b0; 
    assign out[2349] = 1'b0; 
    assign out[2350] = 1'b0; 
    assign out[2351] = 1'b0; 
    assign out[2352] = 1'b0; 
    assign out[2353] = 1'b0; 
    assign out[2354] = 1'b0; 
    assign out[2355] = 1'b0; 
    assign out[2356] = 1'b0; 
    assign out[2357] = 1'b0; 
    assign out[2358] = 1'b0; 
    assign out[2359] = 1'b0; 
    assign out[2360] = 1'b0; 
    assign out[2361] = 1'b0; 
    assign out[2362] = 1'b0; 
    assign out[2363] = 1'b0; 
    assign out[2364] = 1'b0; 
    assign out[2365] = 1'b0; 
    assign out[2366] = 1'b0; 
    assign out[2367] = 1'b0; 
    assign out[2368] = 1'b0; 
    assign out[2369] = 1'b0; 
    assign out[2370] = 1'b0; 
    assign out[2371] = 1'b0; 
    assign out[2372] = 1'b0; 
    assign out[2373] = 1'b0; 
    assign out[2374] = 1'b0; 
    assign out[2375] = 1'b0; 
    assign out[2376] = 1'b0; 
    assign out[2377] = 1'b0; 
    assign out[2378] = 1'b0; 
    assign out[2379] = 1'b0; 
    assign out[2380] = 1'b0; 
    assign out[2381] = 1'b0; 
    assign out[2382] = 1'b0; 
    assign out[2383] = 1'b0; 
    assign out[2384] = 1'b0; 
    assign out[2385] = 1'b0; 
    assign out[2386] = 1'b0; 
    assign out[2387] = 1'b0; 
    assign out[2388] = 1'b0; 
    assign out[2389] = 1'b0; 
    assign out[2390] = 1'b0; 
    assign out[2391] = 1'b0; 
    assign out[2392] = 1'b0; 
    assign out[2393] = 1'b0; 
    assign out[2394] = 1'b0; 
    assign out[2395] = 1'b0; 
    assign out[2396] = 1'b0; 
    assign out[2397] = 1'b0; 
    assign out[2398] = 1'b0; 
    assign out[2399] = 1'b0; 
    assign out[2400] = 1'b0; 
    assign out[2401] = 1'b0; 
    assign out[2402] = 1'b0; 
    assign out[2403] = 1'b0; 
    assign out[2404] = 1'b0; 
    assign out[2405] = 1'b0; 
    assign out[2406] = 1'b0; 
    assign out[2407] = 1'b0; 
    assign out[2408] = 1'b0; 
    assign out[2409] = 1'b0; 
    assign out[2410] = 1'b0; 
    assign out[2411] = 1'b0; 
    assign out[2412] = 1'b0; 
    assign out[2413] = 1'b0; 
    assign out[2414] = 1'b0; 
    assign out[2415] = 1'b0; 
    assign out[2416] = 1'b0; 
    assign out[2417] = 1'b0; 
    assign out[2418] = 1'b0; 
    assign out[2419] = 1'b0; 
    assign out[2420] = 1'b0; 
    assign out[2421] = 1'b0; 
    assign out[2422] = 1'b0; 
    assign out[2423] = 1'b0; 
    assign out[2424] = 1'b0; 
    assign out[2425] = 1'b0; 
    assign out[2426] = 1'b0; 
    assign out[2427] = 1'b0; 
    assign out[2428] = 1'b0; 
    assign out[2429] = 1'b0; 
    assign out[2430] = 1'b0; 
    assign out[2431] = 1'b0; 
    assign out[2432] = 1'b0; 
    assign out[2433] = 1'b0; 
    assign out[2434] = 1'b0; 
    assign out[2435] = 1'b0; 
    assign out[2436] = 1'b0; 
    assign out[2437] = 1'b0; 
    assign out[2438] = 1'b0; 
    assign out[2439] = 1'b0; 
    assign out[2440] = 1'b0; 
    assign out[2441] = 1'b0; 
    assign out[2442] = 1'b0; 
    assign out[2443] = 1'b0; 
    assign out[2444] = 1'b0; 
    assign out[2445] = 1'b0; 
    assign out[2446] = 1'b0; 
    assign out[2447] = 1'b0; 
    assign out[2448] = 1'b0; 
    assign out[2449] = 1'b0; 
    assign out[2450] = 1'b0; 
    assign out[2451] = 1'b0; 
    assign out[2452] = 1'b0; 
    assign out[2453] = 1'b0; 
    assign out[2454] = 1'b0; 
    assign out[2455] = 1'b0; 
    assign out[2456] = 1'b0; 
    assign out[2457] = 1'b0; 
    assign out[2458] = 1'b0; 
    assign out[2459] = 1'b0; 
    assign out[2460] = 1'b0; 
    assign out[2461] = 1'b0; 
    assign out[2462] = 1'b0; 
    assign out[2463] = 1'b0; 
    assign out[2464] = 1'b0; 
    assign out[2465] = 1'b0; 
    assign out[2466] = 1'b0; 
    assign out[2467] = 1'b0; 
    assign out[2468] = 1'b0; 
    assign out[2469] = 1'b0; 
    assign out[2470] = 1'b0; 
    assign out[2471] = 1'b0; 
    assign out[2472] = 1'b0; 
    assign out[2473] = 1'b0; 
    assign out[2474] = 1'b0; 
    assign out[2475] = 1'b0; 
    assign out[2476] = 1'b0; 
    assign out[2477] = 1'b0; 
    assign out[2478] = 1'b0; 
    assign out[2479] = 1'b0; 
    assign out[2480] = 1'b0; 
    assign out[2481] = 1'b0; 
    assign out[2482] = 1'b0; 
    assign out[2483] = 1'b0; 
    assign out[2484] = 1'b0; 
    assign out[2485] = 1'b0; 
    assign out[2486] = 1'b0; 
    assign out[2487] = 1'b0; 
    assign out[2488] = 1'b0; 
    assign out[2489] = 1'b0; 
    assign out[2490] = 1'b0; 
    assign out[2491] = 1'b0; 
    assign out[2492] = 1'b0; 
    assign out[2493] = 1'b0; 
    assign out[2494] = 1'b0; 
    assign out[2495] = 1'b0; 
    assign out[2496] = 1'b0; 
    assign out[2497] = 1'b0; 
    assign out[2498] = 1'b0; 
    assign out[2499] = 1'b0; 
    assign out[2500] = 1'b0; 
    assign out[2501] = 1'b0; 
    assign out[2502] = 1'b0; 
    assign out[2503] = 1'b0; 
    assign out[2504] = 1'b0; 
    assign out[2505] = 1'b0; 
    assign out[2506] = 1'b0; 
    assign out[2507] = 1'b0; 
    assign out[2508] = 1'b0; 
    assign out[2509] = 1'b0; 
    assign out[2510] = 1'b0; 
    assign out[2511] = 1'b0; 
    assign out[2512] = 1'b0; 
    assign out[2513] = 1'b0; 
    assign out[2514] = 1'b0; 
    assign out[2515] = 1'b0; 
    assign out[2516] = 1'b0; 
    assign out[2517] = 1'b0; 
    assign out[2518] = 1'b0; 
    assign out[2519] = 1'b0; 
    assign out[2520] = 1'b0; 
    assign out[2521] = 1'b0; 
    assign out[2522] = 1'b0; 
    assign out[2523] = 1'b0; 
    assign out[2524] = 1'b0; 
    assign out[2525] = 1'b0; 
    assign out[2526] = 1'b0; 
    assign out[2527] = 1'b0; 
    assign out[2528] = 1'b0; 
    assign out[2529] = 1'b0; 
    assign out[2530] = 1'b0; 
    assign out[2531] = 1'b0; 
    assign out[2532] = 1'b0; 
    assign out[2533] = 1'b0; 
    assign out[2534] = 1'b0; 
    assign out[2535] = 1'b0; 
    assign out[2536] = 1'b0; 
    assign out[2537] = 1'b0; 
    assign out[2538] = 1'b0; 
    assign out[2539] = 1'b0; 
    assign out[2540] = 1'b0; 
    assign out[2541] = 1'b0; 
    assign out[2542] = 1'b0; 
    assign out[2543] = 1'b0; 
    assign out[2544] = 1'b0; 
    assign out[2545] = 1'b0; 
    assign out[2546] = 1'b0; 
    assign out[2547] = 1'b0; 
    assign out[2548] = 1'b0; 
    assign out[2549] = 1'b0; 
    assign out[2550] = 1'b0; 
    assign out[2551] = 1'b0; 
    assign out[2552] = 1'b0; 
    assign out[2553] = 1'b0; 
    assign out[2554] = 1'b0; 
    assign out[2555] = 1'b0; 
    assign out[2556] = 1'b0; 
    assign out[2557] = 1'b0; 
    assign out[2558] = 1'b0; 
    assign out[2559] = 1'b0; 
    // Arrange outputs in categories ================================================
    assign categories[1269:0] = out[1269:0];
    // assign categories[126:0] = out[126:0];
    // assign categories[253:127] = out[382:256];
    // assign categories[380:254] = out[638:512];
    // assign categories[507:381] = out[894:768];
    // assign categories[634:508] = out[1150:1024];
    // assign categories[761:635] = out[1406:1280];
    // assign categories[888:762] = out[1662:1536];
    // assign categories[1015:889] = out[1918:1792];
    // assign categories[1142:1016] = out[2174:2048];
    // assign categories[1269:1143] = out[2430:2304];

endmodule
